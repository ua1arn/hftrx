��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�PS&���I�r�`�Ȇ?�O$�F�� �V�i<�q<��tF.����ŵks�=_
���v˷_�a|#�k���[�o�_;��to�_>�bħ��l�Ê&�_[�x�~(c���:Z"_����_lX��Q��0���ۜZe.�n�8=\��d���|����ڸ(W�$^I8�ud¥����*ީ�S^R�_��KR����I��d� 9D�t��O�)��+s��yt5���hm|�l�ָ�I���#s����s$m�C^���T�g�Ƣ���F��p�z)�S���������%\	̉6�@z��v��6�cl����ύ��=Ϟv�֗��Z5<�6'lj�&������frK��q�r=�񖰞��f{���s���r�&7&�9��WXQ-�߇�B�7�.`TMq-|��×��fivp�>lK���헬MN��8�<��9t��M:Ϲ�Y�
59�}d�w��|������!߄�#XZ�.�cZ�@9ԼJ���Y��Y��H�o�+�CI���Q��vK�#p��Y�}���n���Gۅ͒-�=3@uu�e;����.m�OHd|�PέF@�]�a��&�24(�������1��\����ͯD'��<�X�y��\��S'��Ԓ�afc��>x>}�9=p��Ё3'�$�X��i���I�Ԓ�*��u�ޜ�d2��XU�1�7��(�c�0?�	Ǩ�j���.�����K�P�"�&���݄���՛�p6r��o�u��e����h�M3!�����
���;�x��鉴5'�l�_K�kB��Dn�!��M�-��W�C��)��"�ЛM4���F]���ʓ{�����̋*�J�I1os�~��9�jj�;��idfA{���C0�7��'�p��!��?��b��8_2xſm��5���=���&�=���HL]c�v' ������^�&%a��+��?�B�m�S�U�iuN��P���K��p֯�9��4S��U��Oc�!��+T�!ښTFj�2E�8Z,pV�z��,tH8X��ד����7�ǅ�z fg�7͟��,�=&}���M�|"�`ml��0��'�p,��+�5g­�1����&�V/�:i+����d��ۗ� ��Z���D���9	��ޢ�r��8�5�niZ���Y��Hg��;"#vL�\��N��R�q{��'C�1�ǭ~^��!�LXne!��O���h6��>��A1�7r og�;�'�����(-��O�������n��󿙎��5�ȼt�2卨.�7�M���vSSOm6�=	6��/߷�r�����q�&([��?%���~�H�"O���d6("��C��!��<M�%C_�D$w2UX1���\ub��D)�����"���C�(�$��禶�|��-b% C�ބ��t���z7��6)�f����}>I�#�c5��a�����ZLH�qt�#�K�q�p���^`0�z5�0���XT�6c+�?���B�C��3Ӽ���8!H�9/g\�h��3��*�MQ��:ɶ���F��:�c
�H.V7��X�{��:��iZ+4]T� ӷ��p~1���i��G�)�p�WӚ���â-��Z�<�q�)�y�:ێ�;���Gd3u��-Ӕ�{&��B��]$��̅$0+H������K!c��I���pͼr�m1��5��Ӯ"�7�$� �����N�6z8
�F��6�č[崟�[���v����⯫�,Y�����,{�����b��n;l=��6���.�	���^��@{ �>�t��XV�F)XK�����&!5����J&���(��O���cw��/ʻ̈���pk�c���&�:��� �
������Hw���qRs�v��]�t����¯�9�A��WX,�;ّ�f��1rP2ۀ��j��x��� ����"���NEE�ÑӖ[P�\ǉk���Vs�{or	�F��ވ8�6�Q}yn�mE/A����*w��������{#�"�4���!6�#�)�uSة����N��7�R5��ؘ���m��䍜b��a��-żh@�Z�|�PZ�����*��J�Ç����������������p��/b�_ӿW��E 2�=nc��b3t��iI�8 �2������/s6c�2��<j�к9sE(��5 ��֊�=�)BIӂ��T�����܄��|wє��s�S��_��(@��i������^���6�ѫt/�ï޳�*����������g��2y׼�����w�[R"�3����+���G�4ꔃ��=ڳ�LvR��ȸ�V��!�f�}��pj�!|������ĝ�5�Zh����.��΀S�.D��@HD��Ű�w�x�s�sj����R�f���FLe�����aY��@b���Ab]Sd1�K'FZ6n����<��B�>�aPW�*���y�-���L��)�e��ɬ�	C����z�|Crʻ�`G��XY�9�]O��hPxO�PE�E���J�&�JK�\4�B�*�� B%��[�B��&]!f��]!?)pY�œ����'���/�ݟw���ͅ@�	Y}�
h?r�k܃$*y����TDh��4#��O�.�Uq�����佟�cKr��B"�1>�8�,��;����%��=F֧]�K6���OC�}1�mJ*��#B��e/�?͝���� �xk[��=���΢�� �[��A&@ω��2;�(��C����á�d =~��T�����s�{j��y�]?F*�v�a�e(s,��O|��jP���_3��.p���ح�؞��e���K�����>L��PCd������_\�v&�q߉_x���-if���]��T�E��L��w��jcn�XVVBP���y[��߇�j�\��"vE*�����`$a}L��<���d����gg&�5=�ʫ@�b#���~O�N��y芈��a
kE���	8��{����GJ������M(O=*�L3�,B�n����忋v�J��No��,��鲊�New�񅾳t ��^4�#�n�Ҧ֌#���_n��v2�o��r��c^��,�
�3O�gc��,x�G�n�2�ԎΗ<��D?inB��Y����IX�c���aNX�<�]s?�b���n4�jxn�T�8�+��,]��Λ��	��j�8�¡O�W�d�!�����~�D˻��fx�@��+������-��tir]�{݅�`֕�g�rY��0భ�����?S^>C9J�%>jc�;H͐���
`�<�*ݴ�D�����`=����Rf+�hԪ/�r	�
p'��o\_�R�5��t�u�x�2`~AȖ�g�����v��� ���}@l��$���2.��Z�z�Nh���&�(�!3�c����:L��D� Y����͋�S�S�72C����3"uvR"�(�f��B���a�t�<!m��>	C��t�1���P�0��5��,|ٛ�9�פ�
{�>UQd�gݻ��!�� {�#~��C��Ii*�{�z��}/!��	��������c���m�i;d�M8�f�����K�<�)�6ؖɜ���K�VXl���1���6�
�Ah�V��	8���A�=�T��9h|�'l�s!��ٞ�ɮ�U�"��`j�&�dB�OZ^Fh�5��܆Q��)٢(k`f�-�EB��T�n���/��OL�[%sj�5ڞ�L�Խ�����8�B�[��Ef���uhӪ��uo<)����ڑ}�����cLч=. ����U^��~m��`��d�7�u����*1�_�r1��r��T�od��"���1�ϔ�4������`� iLw�Ә5:�;J�����Q�i��ŀ������p2&���f 	��ͫ�ױ}��uf�؁���J	����[�O;�p�A3x��Fr�Z9�DϿ��Pw�o���@17�L�E8 k���j���
}fԱ
��"G��qr���ؒ�ǀa�&h�^Q, Rl��
x(�=����_B������@���o4�C�������黔����O�����C��$c��^�V������x�N�L�$��ێnh�כ�,��j�_�
�Θ��bBg����,f��o<-��O�"�+89�R�$��.բ_�t�R�H%�ƍ�3}UR�2��[t����2t+K��gf|�r[;&Kp�ȫ�.my�PȎ<iEeg��2�l�L
�ոN�X.`�yA8rPL�a`e�ǎ��"����۴jX�ׅJ�oO�pt�r# Zڭ�} f��b�������I���o�_O��[3��U'����EC�p�!&�;�'Г���Ƥ��v49�c'#���$ŏj`� �^���
��>��X'a��'����Z�e�H{l2����"�Lά���L?��9RpR5���C�2�Xp��=<\8&yYI3%�O��/}�_�8�Q˒AqR�L|�td��g@��z{<	zڎ�'M�ع��wx[7}��Gn̬�����������.���)K�o%G�iB6�Hp�ֺ䡌S��0^ע�U���i���^�Z�Y����b�2�h���谘e�F_�|������\�E4�6��d�4'�����d�/���D4�|�`��J���ҏ��Y�
�|�
+�ۈ�F���Zd��Dmi�ϋ+�i6 ����4�ש�;SB���3E�~�I;�Ȕ��X� -nC�#}HU8�q��*�U���2)�r�=�2Oz��]���R����	���et�:�Y�%�w	@d�o��[�5�ϣ��bA��ZGp�)[�	kZ�n3S�z�v�m2�2���f��g���&�it+�N�YhmW�B{�����Bs���ۚQ�l��lbhT�kTh�|P�8�|�f�1F�6j��˫�ƻW �!���2bSx»�W���}/��pG����ؙt��Px�3�����X?�o=����vhs9�a��U=_�l2�+���`�]����5�r����S��^~�KoEԲ��r����ٕ�@�r���(�L�>S��F�?���y/�(�KGO ���a��|��Ռe����&���8:������:���*�l�C��d��{�F�����Zr�P ��N;���D��?��!��t��@��f��)I�>�#����<��W�D��'��D��}D���94��_Z6�:9�~��iU���J��4HUt��,���W���>�7A��F�[���w���R9W�i��1��S���>k8��ve0�יn�T�TQ������l]ݫ����= �{	DJ!7U���O�t8�uKP���p��C@>�iϏ��C͐R��qna�h������xUp-�?�:3���ɿl���=�IoJ�!��K=����qa�t�	�Y��K��6�w9�YU����:Y8�*�ib����H6�&tw����"�P!8\]�[��ʨ0Ɓ:��C(��K��$�B�i�5�jup�dp���,�sP`�&�<����J8�P�J9$����������7�䙁�vrť2��zɒ�^��?�(q�a;1��9(�i�p�;�EI�-��<Ve�̂��<�&})����tw�{�h�NP�&�ϡ-�|W_�_���5rﺙ2��b�bB�(�zn��1�6�9��j����D���d��=�H�b�^���|��H��
���)n����ɳ�Ya����?��n�{��6�c|���V\�P��)0�wMc�gݻ:�U�r�Ă[s?� �JQ@�c%�]�M�9���KMY8Y���!��S:#�0����M~7���>��� 
���6v4e(-�\��9���A�(�tD��s�8��V�k-<��V_��,�N��J2jR�P�Y���`�I�V�9Ѳ��Z�d�C�u� �^.�`�/�:>+g���O���C{�._;\vnU�����5��8/�k|�0b���0�\�K��V�2��^�@R�1��0�:2�b'���H(mX�A%gj^]�/�(��h�vHد)���&��d�~%{ m�_&�����_���N{���c>��������p�C.��vl�V�gs�\��b-Z_���΁R��:�'��j��h�v��b'5��/n�lh"?Ix�W�D�<��m�6�q�Fi�]�:������qU`"�?w]�U�����Ê�P:'��T�3�T����P�rV�-F�.��d�|(�	����
'%��U�R$%\j9K��E8�t�i�����_�B�P�Kii����7�J�K��N��stԢ:&LD���1S�kyjI�C�%��ϥ�i��FM�7_ZVpt�u?�C��n��w����tevG;���8;�Iv�ѽ��~��q"���뼣@��O�jz����]<�������MD�d�1�|w ;��h"}���E��XAMvc���g1���봌�UOH�G�Z�֡�jؾ�0�˕�g3�������3�4�����I!�P�,<�o]��I:'��f?�j/��`i�f�����M"d�_4�
�?���6�i�&�`��TX�/�on��ͨgș9�6q�
������1�=b�8�sT��-��7. &�&u.�C=@��2`�S�[C��R��1?����F�j�4*XW-�(Tk�Gxx�ֺ�GU��`�B֣t	���2z�xo�|s ��q�lO�����D�pYYV���9f
$h�}sY?$������Ro��A��IbY�"ǎWz}�r�<�Z�|�J����K`@�g�)�<pDg\}����_O�!�J��0����Q��2>r����;)b��kaF>m�۠�4�{�KU���TTP��*���x�|X���_�f�� ��np��R}�yk�̩�֘��w�RB���7k�N�@��F(���4�/�Vm;T�I��5�SLX
��^��6���O�qk���M2�j��-b�A�E�񥻙����U����W�T��7\#�>k�f�9ݛ���b�i+��b��O���<�8��<�K�Z��j�a��{�J���{�e�sC/����vw��sp�YҸ��n0|\�iA�s�|�����a$����>�m�}�^ʌ
Q�)�5q�v�ʙb��Apb�q�����T��.��t2_�(w-�� F@�q��l�0=4�a7��Q�`�� |qmG��K,F����?r��rn߾��?�^)ސ!��Y�~*r�ob���,�h^�zq�fsh:�����.��7�fO�"���vZ"S��.Q��8������B �0��T�0Z���q)�#�E(266��ܬ3��|*��[W@&p9�J��(~%Cԫ�?���p�ⷅ�?yK%P�"*�X%���G᱃��*#��k��e¬T�;�y����
s�K�T��������n���HAF[�7�agX��뀾��-= z��5"��P�!-u��=j�B��-�	c���d�c�	�	y�����Kv.�mHr��]�"�Hf��"���Ey9_ ��Y�D�q�W�)W9�՚1�Nc�����=�ݼ��I����1�) }x���,��^���S�~��3�� ��wH]{��;�A�����e��*@I\�`����E��-Yv���*a���礐'�h�o2e�p�eH���s��|W�_��FԴ?6�)9�������{֟ �v�b,Ok6q~�Sշd��pX;r�[���s+����1�'K9�� �e@��?���a��ԅhS8���1��ìS#��_�p�m钰�U6�&��-P�vVzZ�$(�h+�U�٠��/�:˫y,�'�1ǳk_�QB;�>��]�`��s��������{�N�(�{:�5~y�D�F�»2��������^��v�T|7�
KQ�W�p�.`����h���榊E��Ӗ�"�&R{\G��GI�	�LRw-��4�l�����ǋS����d�U1G�����DD��UV��*�v���B�]���\e��O��=PԆ�����=�����u��>=6����[w�9)B���{���"Z�O�>:���6'j��tA#�|���x`���"^K��#��q n���{R�B5�)[�zQ�� Q�{s�����u�]Y�J��y��zz�m��1�L5�0��ᜃ�������
컅��9µt"� ��L/|\�GK|��IK��)nv4�^�Y�a�+�|����y�vPQ���%��0sG�iW����Ҍ�ѯ�|#+W�HQq	����♰\V���N�J	�	�}����E�t/-��Ԁ�������.�?�h,�&B�n��jԺ �
&-�M���V��hjh60aUB�ߊw� ���\�k͙ \��o��GӘ�ISɧ��uW��ٳ��:\���q��S����x
��ٻ�H�p0l��'�k@h��
eML���lJ{b�Q$�!�L��p1���l8��К��H=1C�/Kڮ"��)-���ql����0�@��ɚ�KC%/�)SU�n1LN������3��ڼSy�-�����MT&
EvQ�?Y�zK�ͤ����~�U���ev�e��1���>�Ls6�XY��m�#�L��̖)����i���WM��菉3����W���h���?�{1�/+���#�{'G�)Xӣ���9K�2m���n�/?V���U��IF�x5;�M�`�#�0��l�4�>��Q|l�	�U�_I���}�����NDv(ߍ۝j�#�����?��W��Y`f��$�b-�Zʭ��}�G` �H��� u|��0)�8��[�!�$Kc��wEKu��|������_�ن��w�Q�W"4�E2Hf���g�+Z�U�&$"�*|J8���N���k9v��'�N���*䖋�Kv5ln_�+���N�T�VC�PL���ٍz��c�>�����d��ti��Xd�4���ל6t_�	�4RZud-�vQ��?#ƷZ�&1j"���o(�����ԙ�[��D�=��L̅#
�4&mj�Ռej�GL�w��.��b�����lw�b�d���s<��Kc���TM+�������M��ئ��UC�mI��9��I��p�2H��o�u��jK��f����|U������1���փј�H����"h'���G2Q��2��r��z�T���Yꉸدo���u��A3�f�i�}~f�\�F����O�����~$�Bt�`�Q�vʪ���(�NL8xI:�������%��~ݧ�� tec$� ����p�հ��T���9��^S���}%���d��I��e����0$�<�?�@�-<1}��j]a��g+?�U���l�Z* �]��J@xT֯�Fxղ�,t��r����\<�!s��Żt����r��
��5�$z1RO*��z3�7E���SX���s���S$��ڗ��"DlC饗�H�����3�"�
��}�����-�N��H$	��A1\������˼t��:��SU���*=J���=^�yo���Neu�CO���8ym�ew<��Á�9c~P8ڗY`/�vv��%�)���eYQ{���h
7�E;P*��[��"Z����Y5��
�_+��1��[n���}3Pk�~�=|s��/��9灼��'+&��ϣ�7���]0��������8|�v�����̒���:t��=���Ax�:�	D/�0SA�����$"u��,���-�� ���S8_��i�8mDql��P��`�I�%�r{ĳu�8��C>N�=نpk���=�#�*����u-R.�Q����,�����d�m�r�����<.o�d��H��	C��1��5��^p��,uJt��k�B��_O��Nhp�9Ւ`�vs�FHXN�,��F��<(�&��������Lwu���xWVS��ζ�=ϒm�/�
+ŝ#u��2�E��LRK����b
?c��2 %vӖ���m�U:~�i��r�ˉ٩���a72��D�j�רW���
��.��
6g�Q-�AOv���}h��k&g˒��z��YuǛ>�Us~��T��ӂd�LF
�`Rh�I7~�:֭�ͼRo�#P֋������"���N�)�Ck��W�0��\?.,�I$�ʴP�T.��CѢ������JW�W.[9� ~�}�!K�x���� v����B�nF1��J�w(`r�^���Xt��,4��I��D`��)#
�@��z
pq1�ii`� ��z�#�k=�Vtހ�s���I�����	>i�O�ח����D;M<zƙ�9�����I��������yt�͔y ��XܧB@AZ�[	�p��(�Ⱥ)�y�.L��R���-H�"�˝Ԡ�t�����c�K���\yҏ:��`�e�v��p����D] ��a�|���</$ۡ�^G�s��� ���D���/g����+�TZ!�zY������'_��a5�~��<N_��a��{�h
} ù��;�|��4!���,/�qZ Πv������ޙ�)G�w�����B.��K����?s� 4ºJ��u��p��z�-q��w_��X'��:��(���3u�������%T
��.��Nص�bA�?plp��O{H��|uXk��H����B��5UȞ�P���	�Ư�I9��,d��+�K��x�2��E:-�i���
?��7N�<���5���-	�T �ɴ�%%t�Y'�"��[��z�����hA�G�͚�DhC��4����tQ�����	_��T�`��?ES Iɭj���<�ꇌ_�t��A��1���_ů�SB��-as�)���e2,Z�LPR�Pm	]gX��k?��BZ�eK�kK"aH��w�!�Aܭ��SAy�.����v�>�{)0�%��bk|}I�(�m��E"u�e�<گH�<"x �W@�]�| ���Wj6Hgv؝���@f�H�ąݩ���
�e�s�Բ�G��4���d�����L���\��z��_b*�y��1ߺi�"A��}�����,x��huW6s*Π�tY�%��@�j+Ds%�d�>(+t����3,j&��j���2�V���r�^�Ԅ��WjD�]���#�Q���&�0_�%x	Ԭ�[o��o�'�W4� o�s�z�[�yo��'L�X�����^�mJI�LZ?.�~�c�C�ɭ<30�35h�s�)Uy�J"�o��7�J��S^%���JxB���.�F�H|�@�!����5�3G(�=~U1v������_ŉ�Y�K�(ȁ+y�#�)9b3Ix\���ê�L�ӟ�I<����\��߯6+cwH`��-�۫���8*i��o���c��\]��t|�ldH�<�܈�	7I���aE�hm�k.�G�|����	�$q�f��O�MI�CQ����h(^M��21T�mG��7�Ay���@��x�C�tBc��\�p�W5;jA}�������-IBl����כV�x��Q��_`���p���zc��*Fs'SɅ8(y��l<#���-�K���x�oy�Q�k"� d,Qb������U*�2�$�n�Sl�p�'&<�T�=[;jca�V�|u�.r�� ��Zǅ���"��+��J\�L��Ir�ˈ�����H��$�Y��~}H�T�{��uw����>�2N��]!ߡ|�dX|=h�z	��ɫY���Hh�j	�I§���8z���9�IV�'�9��Z$q�2�?#��YN��dD�}D$n��\,}m\	vo���6�}�"�o��@ҎMH���)kȈ�z�O.�����,?�rn�İ�v�op����/�tt@�Çxf�V�)�$���
��4���	!j�����.| 8���-�&x<��nDCX!�����jV��؛l%k	s~s�����C�r��K��8�J$�������wx��kx��`�B���V$l�s¸YM�N�vL��ݝ��K���_������2�D�V���a�w�^Tܩ-����rwڐ�X��Ea������(��Ǿ����;���z�f��f���HD�OzE�5�~n8�}Y��\�MNK��C2L�Tzг�!Q�g{��ʯN�R���K�h�ۊ���f�i�mr��8&"��V��hI�:R�ί8w� �emdԍIq���B<�f�Ð%�^~��a��
6!�Y�/�e��8�E�Z�;e�;��-kXF_��4:�Tʔ����'2"�����$������j�����Q�6��)Kl_���ؤ�.���ј����u �Ʋ���a�8��Ag������1�ڋ-�g��[&����E�;xV�D�~��L������{���C��n�J8LY,�u�����F���	~��%�&�P,�~��Y>(�3FtQW��7���^puU��pd9�_���V&��Rf�3 �J��Q�L�w�wK��,`{�D���~��@���g�ٌd�@��'��G�5^���3c9���=�����j<;�p)~�B�I���w��G�V�2z�ٚۊ7�o�����>(���-2�>|���Ǔ�n��yD��CNuq>��:E{�������7h���mG���I�����m.kr�-ʳ�씦���.����C��&|�h�5`67�	�)7	b�S�cX'�x*F*��D>�ށ������9ab@�9��sȜ�BQ�X�b.ox�.����mu�t���M���1�P�<ܪ�}�FM��%$�y9��1�/�����mg^�V��;����HC-<Z	�JX=�o`\e�糩��`[\e��O���ϯ�w\�T�n�q����U��.�1���']ߪ�} 6��҉Kd�BaԖ��R�m�[�;�T�7�..^2=�Xo�i�BG�E��E���' z��OSs��3�uOC��>���s ���j��\�n�ߺ�ޙ0E ^e';���h|�����֫Yˎ}j�s�ЍѰ�f�m*1�6�y�rY��^{
����#י�\�;ݰ��~���r�`�$�_�uS
%�5�)�	Ū��򦃁��2Hb�R�7��6C`*+��	��ԑ�[�b
Ǎ����Dϖ�G|gU��Q�?eb�Pc�j�����d}y���N�j�l����˟>8SWS�����w�����[b��p^�J���ݭ.2o�Te:����HԜx~�%jіΣ��$�ʒ���"F�C�NҵfV���[H�{.��E�G���ۗ�Y@wʣ��	�׌cԸ;~D�J�#WR&�����<Ђ�O�G��0@G��TwQ.H��̓�����m�_��Ehy�B�2��u�@uvP�y�HSU9�k.�1:��ѭ���ϝ��@&��qO�I��xv�#X��^��Ȝ�,�Z~P8` SVF�}]W���ap�~�
m:S_]y�e&���(٤i[sk�խDۥ/���4W�Q7�p���E �PH�S\t��恇x>�Hg�rH����f{�`1Ќ}D�X[�>D'�)ګ���9�;�5���} y��'z��5^�2�M ~������&��x"'��8���Z�� [��h��x$�=�f:�>�V�O,Sa7>���q�M_�����z�u��ʮ�^�%�����vhlT���xYF�_����<6Dn�&g�����޼#�K �%p�7}z�;�p��@Dxo���"^��X����ɽܦ��IoČ�
��0f�y\%���2�C���'�0d�D'�}�}�o'��3_�%�ӀAD?�^ะa��iܚ	�O/u�+��A\t�V=~��Kp�4b�k�qWi�W�w/����������}(�HT��V��T�BбZ����o�����~=%)HF�rἺe\�m1���'	[)ZW+x�笖���=�]Pfs�FĻ��NϪBIَ�D��t
��A����9߻ׯj�|���v���@6���\ޫ�64=�Ŕ�0e�*����m!Xі��dR@������"�k�Zٝ7��'u;�>�����)!��q�_�CqDQwㆵW�G�����iD�L�
��rn�Nr�'*x��|�c����� �3�\�[�S��� �j� �@��<y���Jm���h��T�O��FA��w��#�U�Ap�m���NX��#���&���C���!��AXz"+��Xr��B���>OӇ�kM2��lxZi+�� �4ϮE��#èy�m0��%_��lY�;����Q��N�M[�E�Q�+��┛��SF,�r���ٞ|ڧ��e0~���0r����0�Dۻ�_.t�4��4f�p?���NR�-JB͗E��	Tx,�T*���`�1�B����WE�?DѦ�}@�w! �(Kn$r(9��5-u�h�L�z�p��w�N��=����ww�Q҉��}�A��hP�a��1>~.������e�$��q&���u��	'�����~R�]�"�A}3>=����4{!�[��8)e뼣RkEn��X��lU�s��p�հ*�%)�s�t��ɍ��U�u���K����y T�����@�n��7��0m6� C�}��2��ᩲ��Ga��� �ʟ���؁!�"_�Ds���'�i��w�I�B�e�Pפ�2����">�������x�M��;����CK����n�}$^��nh�*�XeF�;��^�Y��fb�A 7��GGedŎ�q�FMQze fޒ�.��n�fj~��+�Q��d)I���FX`��,>)�_�vOXZl6�A�7��z����iO�
,j����7m���U�	�s��qm}T��m��|�+ޣq��!�X|x\�H�L_j�N{٢٣m���ɲ0�iu�x��)w����/�v_��$GVj�I�Gp��f7�Α�,%�e�
s�kϋ읫���J�U`�DO�~�<�M���H�|�N��49�:��l��X��IV��(`��(l/��NZ�)��ex�(�'�/�����=8[�T7��mκ��mxw5&�?��	Q���c���`P���i��ylt"��!��/c,��j��I�u����KRqX�X"Pl��� ��A����e�w�aZ,��0r�[R�c��?�f��d�,�l ��3	k�,-�\a�]Y�$¬�I�r
�I!�vy]H��6��E�X��WZ*�8�=[~��Lj��i2���?�Ǥɂ��+��U~F*�8�ڂ���o�r�Ɏs O�T#�A�B�l���^�!�$�!GN E)�#�:Sr�[m�pf�4�	�@z�6n	bk0$	�L�ɦ~��O]1����㵁�
y��h�NR䆢�ü}��`�鹧�� �X@k�N]hͫB1�6�G�
tf�V2�;�ܸ3�#hOD��R�V�FUY����U�%���L׉�Fl迉����F|���2�:i�9�f=��!�j"*Ee-�%�1�2����$KA�lCc��%���R�ju5��a]��;�����s���-����p�~��_�I3��Zc0ΌzhR
����g��ks1f��.�8�: ھ����c4 z���0� �bS=ɫ��K�9�>_��6[���O��F%�r����y �Q{�Z��r|yh/)�.%n��\v#�z`�*�S i�5P��4����<]��5�]TF��waP����0�K��Nj�����Z���#f0e,�NK=)?��C>s�2�8f�6.����+�h���C�p�|�Y7hM&x�7�7�t�gt�;i��ȯc�~8��7�f#8:J��k��A���c���t0�|�l��P�%ůo�0�䍬��:"�QI��{�Wv,��*����U�J��Zcz��I�]aq��M��B�-7�K_����Gp��@m'F"��6_"K�Hz��t7�qt������ �*���������uG=SF�"6�4�i���ӃE2����S(z���b2X#4�f��乜���%���)y�(�&����w��R�Y���&%��i$jn=�����D��t��q�A�g���[jЧ�������w�3_�0r@��������8A�lD�����ʐ�U+f�7�����n_��#a����+�C���o�k8C��������R����Y)߂�Ch*Ɛb4�kD�ٗ�dc��S6�kv&�~�v-˷T�M��R��9�d�N�w�)����J��k�f<����~Q35i�'��A���o�Z�p�*�܃������#�@��6�6�/ѪG'�/p�~�t���K;��rD~_a 1ñ�[ ;<N�2:���f�����)��3Z`�dtw��J�68�N�g�墵������;3�1�~��`��"��\�9	�A^�t�'�����Q��̳�Um��ޔ{O�)��?琱0�/�DjgV��.�t5�"7'�#�Z���J��7cLH)��WD�G#�Byz�x�Y�k~�c��}���6G`����N�D�5�X�����:1�#˘�8�@�J���#�)���q�Wئ;�xD�4n�����2*^��r���������Zf�&9������΂�������h�g%�d��T�\U�j�Rd���g���wU����H�F��|�%s�]i��@��"�.����E.�H"'�n��N�*UOP�ex?�5s�سP(| ��a�N&7$���j׿�J4��r�|U�G��0*�A7h��U�81���_*d�l��!}�t�n0���zШ�?�
�A\[g�Hɼ���\�o�%�.�̘U_y�._D�2?a�WD��o��h�e�Sr����O�.�r|@�
�[3X�TaI
R�;�W���lTD���FY�3�4&~��䤐�O@����[0�Z���%���h�+KƓWkd�T�VP��|SV ���+MO66�?f5���jC��(�iK��uї�W�-�$F\K7	��V=���� ��Oo���n��
!���5i�j��%v`cvL��@�7i̬��ٰ����G1?\���m^�"Y�B�F��bt�ǛZ�.M�f������/)b�i�(C�&�t�@"\
X��p�@a��B���'�qX�ܫr,�&y�����-�YǺ*(��F�d\�X����3�/p����:�IQ�ŝ3g��	CmM���U�<��$��4�"je�*�|���Y
�_�m��CLd��YƝW�u9�Ϋ�+%���_�y�����GK�'R���(X��y�4Q�A4��� �w�3�]�����˛^��
1#'���3���L�¼[	��x7Rr�HR܂_��UsyPw�J�q�گ�щk�(���\D8��eHM/�S�>�)�I��=������Ĳ��6ہR�3�;�i�:b�i�c�|�&6��c���v�{�ƙ:��ݳ��F K�6��@��ioIt!�F��V�LC^*�����m �_�2d}�R]&'��z8JR�E���R$B�=�p|ݯ��I�� ����	8�9R��C����s���Pc�~�GknX�6��;�[N���� �"��伯�늺Sq�igT�#�H�jM>~�j��}&Mo�n��?Dm;����[шC�2�l(ļ~�a/�x�s|�����s�Q��'�*�F0/<I���K����aע}����e��l2e���IC���3ז"�T�bҵ�K��?}QX+�/�z*�X�0�ך������~�Ѷ=<�	�a��U������_��N�8�w;��K� �Shȴ̱ͤ���̮���N&_��r��h��t#�ݚ�Ԛ^I����H,6��3b͕�֩��J��*d��_A�f�;���W@�k+�l'\�t=��oE�=\8�>�|J�1�C����犐�֦����7ǂ��=C��!!�sE BHkC���O����:�)Ē�UNBr�
ܫ!⎔I;s>=ڣ]�k
@UX	�1~=Y�h�	wA^tċ&�(ifpY�}l�zC��'���P2��E��R����ї��Sp�5!(�����gGUsގ��/IP_9�~Z�����m,G�KV���4�Cl~�d��%%Fa٨�(Z-̏�!�곹�������tt�V�G=�G���H�(�x���c�'�$�n	���N����)�{Eh
�,���*Ё�.�Ъ@�%��/��Rbj�t�h8��W�Gc9#.T��VUf��<��~�fjq���*�ʥ� 5&pJP��-G-y6en=4]��:6d^S��̾Ab��_����Ȟ�%�"�D���ǻ"��e�`H~�W`�����W�u���n��f�Rn<���v�GKm}M9�4}�]���D&h�\	���AVjm��@��c��7����$�����oaf[;1#&�=�w�y]gF��W�"���0z�]��6�^j�j�=�y;$�?m�W\�7зI�K��t?��i2ȷ�;Bf��)�_�F�x@�����8 �;b*�wE�������.�e�{.��ؕh?�e�]BF�$0 ��K�����E�f;pB�M����y{��7�ÇH4���}/�
�Z�2g24�'ӫF{�2>Z�#:q�w�[���׿>w�S(� �ǆY�YO#��
�Eᩉ�?9cr�kN9|A��&�)���1z��Brw�Oj���ui�3� %w�� �F��An���e�k����7�]��%-�6V"��eR��{���,���Y�tq`��Y���[N�H�����Ϥk�oO�c�{��"� 2��P����,@k�u4�R^�*�QsҜL���I������a��e�z�Mh��,\��sde���XK9��ķ�
omG���4�襸��:i5�'4F&�IJ9���B&UȾ�i��t� ���;�(�}����*��\
j㰜�Y�Ya�fo�ι��]a8�����x���R��o#�i�4�@�1�b�U�t�Գo`Ƒ�3��v�����.�?=,tx��s5`�鷘�1��ײɪ1yz{i��Z}W�^�
�O�A��B��*,����7c��3aͧo��2�rZF1��hV�Nm��}]�V5��%�+۳c]����<�q��Ĉ���#�l���e��Z��d�G�ӓZ,�Z57˳��i}��%)srsG�����y�9�O�� �"�?$y����s9*��>�I�mlx������m3����(m^a"��Yz��(����o�RR
`f�d��!���ǩO{j��}�2^B�5蒇�����t�G@`�����;��АsRF`�e�K(Q2A�q���8T�s�<�V�Ӕ��^�\"�1z*}A��j͝�"�8�koՀ�}ڴU��b빭�� �`�@̰�R_v/`���f�M��Ru2Kh�	��G �|��@������I68�k�%���S6�(�O��'5"��H"ks����<����uw�?��UK��sg���<U�F4�.���L$��q��UF��'���'�d*C�������������<��6v��֠���8�,;���=x�Ê����雲Zv��PC��J��N�P��8�ɡ�䂩*.kbq��?hs��&"��̌��A���z�� �R��;�*��n�<�L����2���K^�w����~�e�{�;׷������͚+^x�-|����.cR`DڧF�_�V�bZ0���)>���?=�K���g٥V}����n� �?wk��5r�MđIrY[�ȽP啯%{:9�7P:����O�U�a]�2d�$���r--�]t�H���Iʩ�n�}�p}(�#�<�&�*y�Ohj2�H���u���y��,7�B�����%��֭S�"�1�[��t�����P�J����a�8w���i�G�p�\E֊��VT�F|R���|ǻ'#Q�5�
s�M�xu�gIa�<��V�����1�|t!�y���btJ���pï�5>��8�����y��8��!�ViL#Ƕ�7���D�A��1�t���JQ�\�pZ(o�?�5�ìr��g��2��m�%e��(��R��띵G��/��G���h1v���!�?*D謟��
ԋR�$�-`\��g���[�&�m`-�a���N�;�2�E������^_�ծ]�
j��Q>��#����S�x:�В���n�_��4���R�u[��dҗ�σ����VT(F6x���Bi���!���2g�`��p�;*Sq�M��|���u�~���wƔ�z�2n�5x��AB/�n�k~ ���Ʊ�K*���ț�9��{F�P٪3���.J0�B�W��v��ա;��JD�a�����:�<�+c°b��@��95�;s� uݙzP���6	�s*�s3-��Zm�Z�x>7#rg+5 �K!����?����t'�L?~��^��MeVrO��6�%L�y;y�b�f�_���<X��=}����Q��_������Y.�u�c���\+����m�1b�S�p5N��06��a�߬q'3�aeV'�r<�Wׂg@��8����|������P7�~�;�{)��#|�2(|��Kp�|U�����-3d2#j��҇SQ<+���F zX�Vk�����*�F�P�.�ҥe��MZ@=��k[�FXX%��9�n�wTbE�3o�Y'�gBj)�sC�Br�Wbk�P���
·��ŋD�C#��������
��7u�{���Wx1o��Kh�NN��Ns�98�I��Y{$�t�6��M�EBD�4�ȏ�q�'^��"�a�����9���,kn5� ����"'�ZWa�ؿk]:��El��G?�sN���:���`�1N�t19d�e�²W����+�Z� k.�S��~�o^�H6�BQ[el��		��*>5֕��?]��5>ώ5_�k�iS$蒡�tj���A�&���*! qd�n�:��547�ݛO���+4�� $�F�!	M�#�)O�|�'̲�;��mpS)���� e_����gp���ʐ��r���6��~&�[�(@,�Ƿ�DБS�ʃ��4
w%���׌��o�赵��;��Fȧ�	zv|��<�Zb�d�h)���*���䅒