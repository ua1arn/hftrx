��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�#!��{(�N[V��/2:DY��6���T�'��:;�5(8���$��Eʀ%���4e�p�;��a����^JN��Z0����> ����Z�� ���1���C���Ղ���Z⥃^��մ��%���ݎ���
E~�(6���B���$�i�D��%����?f�G���Cy�����J���ǩ��5���z��d�޹��L�t���M���TD��Z��oW�����l�$�+{J�M〮�
�qH�37�t��KN�s�$D�^��E�޵�Bl |$�[�Hʽ�y^I'V7Qt'��ѣ|DA���Im9�-���Ww�qG��>�soҐ*��^h����[��<�Npz�沙�����@�-���\(�fR�i��rDz)�J�}���Tw�ǳ�u��%��	�w(�U\���Z����u���%���9&�c��h��h em��N�(� |���i�L��t�4��b_���A��7�VR��Vr��R=�f��8�%=� ���)6Gu@[��i��U#�ޔ�-OS��Ӊ�v8�'�w�l.7�ʋP<�k�<"W���	2��X˵��
2��0¨��q��	Ы{�P��m�	���%��K�O����[3�;c��D�Q�I�PQ5��,��ձ�{Pb�#����3���51�Պ��EAyl�������xZ��⑞־.x0����[�g�٨=b|���j�|O�<�]��tԠ%��h�����>l$�'RG�a'g�ա�����������N�T�s����a�
�Ȱ�e��Ӳ�����D�9Խ]��}��~�5�p� �U�s/�i�$AW@-5nMĨ�U�P|���Rs�
��k�`%�"o�(�汢�ߎ?ի���tDg�*��3�f��h<9 �,���d�v�0I�KWI���B�(W���[jC�^��b8V;�ů\fAG*���{���fu�Y�$�s�z����$�i\���@�C0��z�@b�	�`�4a��c���%I��a�r�_�v��?���S�H@P�H��ݕ	�y�8�]�O�T*x�x��u�hq�D�l�X���g. �f��!�#��2�V�W���b�L�>��A�V2d�OI�U|��=�$��Mx�/ӳ�^����S�ꘆl@&<ݚ��պ��`9�cۍk{r�%J���!�܉+ۢ6�.Kw�d�(��^i�u-\�5s�v��u2���)?U�}LB�J�x��øc��ߓG�@J$�>�q�9�nX���Q'rP��q�ZP�mF���X2��Q�v��9+����N��&�7�H����sw�nK�mS��
4��·�ܫ���'��H��E��G�w�T~�eRg\��u��`�@���e9�,�Z��^���p����ލ0������T���gG��k:�����˷���1�����&眰ҴhH�(�����q�傼���r@�$��@����M�-&�s{���Y�������6�퐖��=T�����/���+�S��k��>�g����m��j��;��"/�T*+��8�[�㫣SvwVXkn(!��}<�5x��0EȜ����q��b���kQ��t���Z��3�;�1���A}�=��f�syu�R�֯�%��C1�ɣ�+ϯa�e[���D2�4�֤��v���I3����G��G�@e���ߒ�u�ܽ�&�Čӗ�w7���#�쑉�Z�1���ׄ9�> ���}�:hk ��p�Q��_�0R��cVJ�;k�CŊ����J��4���n��R.�'�<I�Ǌ��+f��h�����$�¥n��ȣi��x
�ړ���\lu=ZK�JV�,JN����ҕy��� �^](���#�U^�����~��{����	�΀f2����vE���jL?��d�ȵ�nXξ�Dn��}��K�E봽�k�9�7��vʒW%%Ki��||����r�j�H��=1�s�T,�������pA��:�s�_�<`�w��]IC��d��V�U��h\�� QЭάc����8)*\���I��F��=`	�tǱds�b?l�R:�O���%n���^՛���U�+�hĔ׵)�;���DDn�Z��O�%�[�Մ/�]�]Pq7�>4����j���R�Hs8��@!	pBE|Ll՗��/��VEa��$Z��J I�X�ͅ��°Y�<�2�5�y?�*p�ZW�Mfk��r����ہ�-�����u3��es��^��1��~-��'t����HQ�]�b<B��o;��5Y8A���-��:�^Vo\���U튒zѫ�B��(@��2e#�b��V��a%�2��B��ƥL�o���Dp+#�{QAf���S�c����t� v�ֻG��L�]�~0x��J;R����a,Л�n��T2���I[�M��ajP�Tg�Z���*�@(1�Sf�MP����vp�"�j��5|jb^��pMtDB#ǫ;Co�u"�:ӟ.��w�V����Py���>w�
Sm�tt��y�(�I��Q�~B��A�=1��q��꙾bK۴ 5l�v(k-0�#1����1C����kE��cm�b]�Z�a�̱9����}����]=幘+9���G�D}]�8c.9[���ua0w�Q��T�*��{�i�>�k�0Aq�MqNx�� ��ka�yE;��oŽm�
6O��P[���ש5�tI�����-]�j-�m��O��w2�t).����9Ɣ}�f����mb����"	�pr�����?�n�4���0��k}���/p�������Dy�6�nL�)G��ץx�����r�+�_6��.U�h����E�swp���#���C凓R]Vd8�ǣ��妉E���D:pi��J�8Ov2�U� 3�ܸ�B��
9���s�޷�.Ke�3N���Ȋ{øNo�.���m�&���8��6�̤R�7�.�x���+�̉�+��vnҍ�q��;�@�f�c�|���wJ+��gg|�n�x��z���}�t�;k����7�����I��j�>�}������V�\��`ם��.#0m��D���(��$I�`i�I��KS�Yvf�>�ρޅ�8��O�>�%/�B7������+_m�(�w�eC��)٤`t���[���7�BP{���.�m'��8��|�8�����܇�P�<$�u+_�N���.��E�� �T�هd)V1:vsdn�*- BO2�f���
����r?#�%<������}?\-����l�������7�j��=�_�����'x�Λ5ȡzH}�b��gi|�޹��C>T�z�顁#�_ia�w���H���� � {du�h��_��H��R��Ҏ��n��[]Ml�X�$%񭔈"d�Yr%4e�U����Ň9��}G6�i�``���d&��n�fO~�*d*&�x�z�*��� ��d�DaH{w*E��0����4��V��r�4c�OɓB���L����4$��K�����f�[�[��I�TP��zrAV&k�L��%N�t*>�{F>�縔lQ$hh����F%Į��u`9�е��>m�Q�P(D���	@�#|�<!��)s�vr'�J�[>�}H��Ms��⵪�j�B�]�:C-�p�O�q�'E�B�G����H����V�;S1�#l[��P�$�|��N.�64_����^�U$JSG<ڝj�6�
��c�����Ԑq�C5�&�����<��mKk>��=���U�L�����K�	���R�2��h]ia��:S�ސ})/-���u��ߑ�~���'ͥLH�������:�!��|��l`z��K�Vh���c'H�(���Vm�6�0��_5�:Hi�YuU����Y��^M=��Y�z+��@
k�pn�I�����;��eĚ{Q�O�?����y�ø�����6<����8��=�$]<$�}��z�%	<]w�:,��?]33)�<	�h� �-]f��ko)�)�dq�V��΀��?���;B�fs�#�߹��F,��U5�����1�.��t*Luf1�F:'�_D2��N���æ�]Ӄ�l��������7�"��5�(�~!w�l�^�wrǌ-��i�������s�ȯ�A��C�y���֍�����	�hA�a>�CQ>X%�<��d���z��mhsC�owm�d�nE$�������`����}ŊQ6�]C�i)��ɕ�g2N�Q�aݟ1!ᠦB%�|8"Α���&!��
Tp�d�z�׹���3���C�-��$�9�j�:G:$�n�z<E��pm�M�;�J��i7�
��5�h�箍�Qѷs�Ų ch<wi��F���H�ڥd�G��שw�Rؼ}�WS+u��Y��ix32��|�s�B��v��Μw]~K��^����`��[-έ]1B�, ���^�ZK�f�\9�7��EJ-��V�c�К�@ۊ˒�, �H�$��`����ǲ#F����۪�~R4�JW9p5Y����8��Cv���&�����L���/��^뻟�ݟX~h�d}���Ak&LC��;[l�؏����o?��p���O���:��/x}u䍝Ь�Q{,
"}+�`3{�^G�y�머w����Ń�����:�9��/
�>�#?W���wթM�;���k*tb��!@�1��׷���(	M Y,����= '�]��¨˅Xʂ׳�^7Y7��j��֤���`�-��km���l|���n�(I�mU���/��S�����fF$�Y�!�I�����`HfS�ǵ�g@��y�x
iS�ˈE�PdU*К�r�\����R��cv�ͺT$�#u8j��h�l���`����K��砆G�p�,is%t��Y��g.�Ͼ�Wl .=��]� e�[�`��q�ܐ�J�)#�ӷE�5��)�׀����[Zʻs�;�=�Z�M��;�����,$���:$�	@�M5���Z\Ϛi�Ͳ!>���f\��?#���c�՚��㨀��@]a�l<U�`�5�t"��#
0���dy�s}�"��Lz|.Ϟ��\�LL��7��Z������Idv�-W����"��;���i+�!&�y<`c"#�k�L�n��9&P�
j��+z�=$�~������PP��#r+I�uP�u1�f9v���]�+V#��c�� !b7��`��<?�Qa�9�|<;c�t��%[=�pJh�k�����A�HJ���X�JLv3E���
��e{���!��Ҿ�_Ts��D�+/���VgD���El�n�`7����(�8j~Э*�1ez�zM�'�?��4U��Q��F]Ȣ�beC+�-����(&>�p�u�����d�>�[OSXm��*�MT3�P慯)\�S���>�Ӧ1����$ +[��WC푬�Mp���PO��ms�4*՜ٟ�Pk�5����8�L}A�$71���UP��+ '(���v���z��-T�}��)L�jPp��kQ���wY���~͸&$�S�ߠ@��*�J��N�^���Ӕ��0�jݥ� ��-�z���`}�CM�[�.ag48��N�:�E��l����t3A�}]�T���!3�8�ΝV� �Q`��&n�n���z��h�u�Aj�C�gY������1#�R�K��7{OO�M���f��$;�0�\�av��[9pM���w�C�G��^�A_[6˔o�x�l�b��k�!�7:>�����А��w��b#�l�r�3�;�`��<)m	��?l��a��_������N�����#���2oI�󥉚����%��s2-ۓEr�o_����Txp�.��_�y>�������Tc��Lt�=Y ~p��G#�"��
y"��d6��ߞgDSUL½�KR�-::��B:�X$-�t�8Z���]��=����	Y��-�������EтN�zUnW���n<A�a&��^�x��'����<�\'q2yr��/���}h�9����>�#����1���[$�%|���"vyw7��k��D`h���M�"�҇�����˦���]H���е\y�x'������I��� �1Q�<�
�xO�����9���x5��a�c�}�3�z��H��0����}���\�q�;��tn!a˛�G�`T����>�=y�d�Q,��}~!����KẐ�]{I<���s������'���mF�<�ʝPq0�Rg*"��'��M��k�ŕs{^&��h�ha����u��n���������23�=�V����l�"z3�� ���?Je��+�a2)tD4.h*��-L��+ɷ��r�/ʆ��*�¬����GQ�f!|��0��C3���lƠ�䲛)''l����HSV�'
))K��D�,��kp>56���IH~������X׮ �+[/M�1���b~S���7;��--�.���(��fX|��8h���5�@`Q���+�%��N��' ���U�f��4o��eH�}�J�y��Ć(�W�mB@��,��V����0��y�&�$'ߧ|4��U'����@!�=�h'�O�d����}��%�)�X�����C�E��W�J.Gz*��k�NcR��
�`z�lRw�gĎ)���"�׳b�k��擁�����U�l9��"gۻ���KQ�1f[�c^�v��t3뛹�v_L�6��L�{��>�m��W��D�5�@J�`���^m,��ݰK��*HE�m[�7�T��,�$Ɏ�P'׈�7���9-5ү́���"�j�c�����P�,6@0xc�lW�пȕL�+κ�haA������%T��#�d*�?yxyooBX�9�����M�(M��U���Œ��
�8�]h�z᫝�)���u��{?��4.Gl;��gR<��J��3��{e��(;?��cvГs45� ���t���-n�q'��O\�G¶я~t]d/q��U6��S7���]��(5�J�}#K�e��$q�"s@�/����K���ˮx��/7.nD"0C1��ӊ�dC��Y$�v�W-������â��~gL�?�=����PI����%;�o�oN�25wa]�B8K���p��(�n�X�
���w	�-QB�衛�&�ˊ�� ����K�f���bƜ&f�ȩsJ���� ��߃Ж��=����D4��a�C�b�6ˊ�ƨj�Dl��ku�I&�	�`V*H�{([�iT�
��G#'�5zQ[����$E��6]�R����ն��Q��J��ڒ!͜���ƚr���3���g��]���ᡄ�ԸJ>׻|���0e�}�k��6&���kc`��