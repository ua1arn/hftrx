��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&���������})��l^(S,�]ql��;֡'��m�F)��T��i�gkXc�4q~�VWt���7j�9;r��W8m4��I8�b�)�Yc��e����G'�ғ�d�H�4c�����<�+�%M�%�����I�6�}��x8U�>�ȧl?�,}(��n�1.X����RFئ�)6�����e�X��1�h T��Ӕ��S��-�R�HYp���:9r���0v�s7���%�2f_���	���J��Wh��O�>�
v�EMK�bGlGQ��$2�{k�)�0y��)�@ �u�x�5Q��ʀ�����A��֫������실L#Ӣ����e�G��걔v�H��Ȱ�7�:3R���S<�����3��sV�0} �x�v��S����>�q�SG�U��>�Hh��?�maO@�Թ�2s�l��r�����gh���#�H�jHM���Z"8�v	�j�`�/�k
����X,���{J3�,�}Z� �r�j�7cMu�����;T����tg�=��N%�R�Fw�r�~I�錇��3�K��J,��!�}�j ��%h�5�?	���0��~SEH/��b����w��Xch�����#�e�n�袳+�1�T�{y,�HA�/iMs��R�zR%o�b���}�����W�����	�/2�.x���m^6<�'(5T��b@��A��W���$�hZ�2��b��AY�Y���a�.�9��/2��!1Kg�P���p�Q�*�7�2�&3�(�����MAe�V����w�;�w���ן����W��D�vi�HP73N}�����@j�z}��-a]��Mhbd���;�GԊO��@)o;�1�Oy�ũ���s-���J�N �#����u���ً/2��xF�k3�M(�xB���6Kz��3*�"d��9y#~#p�I� ˞GԺ�ԡ�_ry�	J���b�<�/��UH���>��\D)@��=�C�k��%������N�y ��b��fc�/��b�8��O�y K�X啈,�����p�	���_-�6.����q�xp+6o͂H�7˽7������h��u�0 j���T�"_�p��Z}�{
-��I�J_D�-tɈ�zc��������(:)[����sx��:NW���ǧ�!a��?����U|���8��n-������=^�z��_CVfZLsZ�����'H�s�ȼ&�7����fP��9��6�� ��ҩ}����BG/%'Ѯ�N��,�z6�P�8B��;x��ș��!�(�"�p�,�y T��𒾚���=���*N�/$��7j��7�RAσ[�N��4�c���~�q�ln��0�����2��mH�l��?�]�0�!��ܯ-�na2���x���L���e&1�l�ńt��nw��� �KX��E���sP>/�杤��U;�db�=���=H,�YNِ V�w�uL�y����s�U�lz��gS��s�����sz�C:���VۯS�GmA��p�H]�w��0)CCY��^���m4������|���-q�6�u8��?�Y!�B�����/�S��Y����tbT�QΘ����g/-�����,���R�l�ęt��N"��E�;1e,2�P�5�'d�z+e�G-o�|���n�vu��T��.���{狉�~v�x��%?ȥ)ǆ��6@����F�Z�~��w���C%8tzɱ��@W#d�E�$n�{� FA}k��^V��Y�j�?�s����~�!͑�:]�5�����ֿ�J��}r���yN��ÒWbOo�pEr4�t]�8�����=]�����B�«ڜ�3���"���ę#�d���(��p�ŀj��
ѩ��܍�7��������N�cI��um�>@`���`������>>ɯ�P��MS
�+
KS�@B�|fw�5�����C�����q��v��2�'������b �#w���(��*B�
=R�Qg4z,$�_��ï�!\8�G֏��{F�U�p���Z|�+�
gϠ�6�� �ۤ����@���ܓ�g�:��}���dDOLA�?�S�"Gt�@y��b�b�݉�*���
�l�L��u�g�*_�G,Ǣ�d�-�u�yC��(���?�3y�@f^�ʓh!�vZ,���5	O+�C��	�G�[�gO�E)E1 I78u�|���x�t���dփ���F8��Ɋ�kw����h���ؗ���<����%-�7
3ԭ��d%�}L�_ԃ�f�m�)��?��� j�7��aT��Ym���:������Q��<ӳW5Ǜʮ�u,Kt[�*��*e>19�EŘ�������=a��d������]��q�mF���C���A�I��W�� &�����~v�j/w?�� ��Q��Z0����$���� �a$oKu״J9��8[b��r+�,q���P%���X�]���L����N��<ڄS�η&�M3<�t�O-~Kh�b����Y�RX�4�����?݂����4}r?~V���dh,j�sJA����%�d/�;=�K�{8>F��N�q��eB��y���� o��v�1�#uf��_2����D��F���x���`t�)P�οK}I]�;�܊�#ɟ��9�7�̓B0����HY@ʷg���p�N>�Z��D���A7�1߬�:A��|Wǒ�k��t]{^�8'�K�f>�aݐ��KI�Ɛ�ٲJ��Rk��0�P=�JDh����[A���͘�!>'1��!m�j�t1Ӂ�,%�ry�c�U���.�0ļ�t ��S���P���eÝI`y�j�'?Ԏ�+r�,�M}S�ryyt���ʶ�<��l��������9�M�xpY���/{��v��Ӎ���}��\B�ίoG�4���\��́i��>o����C�o���^�� A�u�cm�V��v����q��]3#,��J��\:"�R���L�>R�VN���2Hcln��QG�щ�pג���EV�.�[�tq�`o��J2H�43��^�P�)�~]h���w���eP��39�RS����eJP��f�I!��B�n��l�����qZ)T�,w�65�Tb4o���;t�M���	��`?W�	�(��:���\FSc97[���d%#����L�|������r� 
.��o�/�&��:i}q̻�ʗ7ۜ�Y���e��5R�1V4���"'��1���>/�y�v�����RF�.׽�4l�����k@�~*����]�$p����2�����<s���D�d�p�	�L}�[_�j$�d������=K�������!��#M_hj^��F{���e��W;�V\����UDC���@<7Ȧ]�"���т�n�2f�\�+L�&���(��7�s;s��C�r6D��i/�rNF��
���_�ė�4.�S�[H�D��WĻ�[�p��@��:��k��\oO \ R��C\}]h�4Z�=/����0���F|/�D=�?�+�'!hE��������8�'z����z�,���ɥ$�u�݉L�]���Jн�j� h�gN�+L6�*)�`�4SP�����k�7/sF���Or9�m7&T�A::�Ä�s߼��^!��� �JY�h�Ѹ%�R�빩x�}
��>c_�?�Y��tf�}Fx���l��Yr���w+#�nh6hK�&��I������w>������w�M�[M�m�s�UF���Y�U,M@&o�q�=�O����,r�<nl���㞈8Q�.�C�������i0�d�2N�I'2��Hv��V���^޷�	z���~y$�T;���?�ߐ�3��՜c��rc���/��p"U�\⎾lW=�'^(l��ل���]/z̈��2�7/���Qm_i*T�Q�{��ч���rW-��|
y	��~r�G������śH5˶.ڂO��O��2+,����`fCAw���=�_���3>��K{\���R����ȃ�c��B!�g�8�o��։���Z�U��D�p!뙪��4� ���ͼ�y"�e�u�F9e�Q�`� ������N���h�M���%'�A=������H�	�f�p�k��1���E���۟���jfd5�D��"�ݧ�{���|:�G�Z#$%�6�l�F߷k+�F���ɵ���B����00,��M>D���+q|�g����8�h��8��1��z,e�q����oP��{�@���ohs�t�%���ԃ;6�HG�u8N�SO����r3� ���ɿ��pD�ߪ��D�ZD���*C�V^
ժ%C3��sJ!L����P��.j�G@'N�:zh���_<k��P�ejqF���,`]P�}i���I�������Yf��%�@��������h5݅�J|���Կg��)S/�n�4Z5�c����P�ԥ�-��M9�b���V{�N_���c����݊&��=�p��DB��9v���,���8/4n{��ͬ%�h�!�KT��ML�p�,�V�3�`�r׼fI�\�[w�ܛ��W��]�����/6Uq�1���8��hj��^u�����Q�(Y�Ƶ��ZĲx?)��y5܈�:�3n'⸐~Iyy�4d��UΥ�U4u$�ո��q�RDLZ�ǧ<x���<�!��yiZo����:0P�]�b�K�Q�9k�����=��EA-+�.��f*�N���W����#}�y1��������!G���f���7�`��J�֜�~��Y ^Z��!�Š{���i�g :{l��o�]�������#ª3���_��PY�n�D�C�a�'S�c����D1���嚂������j�gUJ�Gu�)�(w����+GŪ�c<���~EJ��=�1�`��B�t�0�K#W���mID�/Ab.��V�e
ܘ2�1����&!1�ɀ,&�������,���Ee��֝^�:�=�S��Q�M��F c�{�"�6CBvh�f����լ�� z��J�Ϫ��bqAr>u'��B�>��u�m�Tʁ�c9*���Ӹ���4^g�j�.�� QH8��or���|��].�m1$0��z�&������F���|k�M����I�cha��QB�Lѷ��χI�k+�n� �?�7ƛ_�����l�,D�8��d3� O���WE1ZNg��GeQ���Ń��XI�q�4�FrT��X6C�_'�Bͭ�������Vӽ����kG�Tџ����nǉ��T&h�LZr��T��͒��[�EV�z���!�c�wB#/��Ј�Mk�4��ЁJV��y
.*e�9�['"�̔���<�el�v�w#ݵ��Զ;8��)�u&�Q���u�]p���1d��|�Sp��<������+ڸ�	 1���E���N�X����t�Ѽ�l����%wS|�"6��ʋۇ]��p 7�D8F�b���V6\t��:U�Lp@U��P��f�0H":���/>�ҰR��$i�����Y�.۰Tr��O�W�۫�?U;{+rd�!��S��t�IB�`��^&mNl8b�u��\u��wN�9�6:.'FWO�6�W�I�עI�h/t4d�,v�`�;LV��Mgp����ɨ�$!?��!o�T5�)�\����/���56�I�=� ��w�(��d7=���q�\�$7�=�i��6�?�ԓ����j9[C%.I�f�����$}`�=��I Cx�������ؽ���rK�<� ���}�3G��v�M���j��,�d�����D<� lZMק۳!�Y�[�$�T<}��)�݆��u~���cR���+d5$N�
���X���FA��ͥCb��od�Ҝv�Z�Ƃ�!���Ҡ1+�J�/D�]6����"1�8�^Rq�'*�I˱ok�ad�o���tZ��9��|�b'��=���@sP����99��ш�����ݟq0�bd��!��?&���S��\�7,M}LO��Ѡ�խ�#�8N�z$��|z
g
�E JBEA�)Y'�G;���~�nʁO�uzvc<�sy�|X���S��v�c@��_t�#���VȒ}�p�*��d�r5��o�0�G��Zl�k���-Ǵ�̦lv[3��̀<Gl+��<���-'`�٬絪��o��n4xE���CPjI�~9Oq�?y�t$W��>*��n��pY�Xh/����[����^WuQ��sH|Sʥ�O�nmcP<���˸ٕ����]Tb������Sj����)i�T��v[^ �>�\sJ$�N�爡���f
�T��������b#̦&�[�u�[6&���c�E,�������X�Q	Ǳp�)����v+EQُ̋�?��Щ���O��'d���V�p����I��G1����x�����Z�oI	�N7=�!��7%Q��5�*��@�,=���T�mu;DK��+�1�׈�{��Q*�� Q\��H|�!eQ��P+x�k�NW�q���C>r�����ߗJ*e��3"t�%3�pj��hW����:rU�-�O���jy�1�t2b���HRK��fgT��^h���/���zJ'����r�w�w�ٛ�譀h9`�ױ��A�����a;����;-1�J6~���:�H.�����nX��=B�V,�?(�+�
��4�@�+�8"|$��=vZ*�1��I�7�4ן�����	��
��.� ~�6,N}3H��Zm��?��&' C]�|�B�)�-�1���80sٗWo4���`\Z��t�ZW$̬�]���l�p�=�����4���{c��&%0����	���Z����B�[:Fު���FA�8���܄�m�6[��C׾�|}"rL�YX�C2��I�����i�;yp]�6���?%/�hW�������
����S�Kÿ:2C����=|�@�C,�V�>�₊Ԧ��[G���K��K�L5�,/�B�bE2����$�E���h�a�K���J=��X����U�墱Z�~@�O��x]����w
 '��'�+����X,�S?q��}���������:��#?_[ߕʆ�R�}�6?�?6�{Ü]�q��%�HG]��/�d`Gj1j�Y�R%5iI�= 8�r ��5�_�����{Zi���sw�����,�k*��=�xr>���&�ch,Ж�p#Ҭ�G90O�};
�d��}��K��?L👧^���v�k �F'��?��&���Kk�{*ŗyPq/��k��#z8��e����1~Q�fzስ�H]-N�i1R낻eK�ӑ�2տ7���{��8:�#���$�6�S9�
���m!3����$L�ӕ��U�ez-h���D�c5���YNL޴�i��&�˰lfbXC�*�꩖�ϡ1r��G����dҜi���C����u=�Õ/�z�]�š��hU`h��4�'�s-���&�
MW}����Ye��N�5�����c4���r���R���G�@��n�uދ����$�8��D�,ch���t��hZ�a�-��ٵ������SB^�,	B�0�.�5��[�<�?PͶ����+K�N0������ߛ��z���2a��2���OK�4]�PR�G�yj���ِ��_��	)z���\>qܕ�(wC�`�=_3�(���Йf�y �pp��!�R;@��ԲNZ�������5��0-�r0����^��� ������@Tu�o�����g.�M_���g�&u��hr���i͓/e�ư;7k��N�ۚ+eO��iAQE0����ϓ�{~�ȕ��",Ԝ%v�x<�FJPq�J�V`�<�yt�X���+MK�L;!Q��ݓx;����ls4�E�	�7��_�NЪwn2��HY����2�|=	��Ez<�rfA�a��Xix�V�,[	�A��/n6��[��2�+j�3����W��Ok"کq�����9�#RUg'i���J`Uӫm\l	ڲE��$+v��(�E$�fޞ���k�?1�7Mʹ��������O/����/�u�IÅ�C
0�t5�a1��,o���d) ��n�{��D�t����{%�R��D��t����I�D�U"y�ȹ#P��`��>:u�	鷡0j�Y=}�a�`=�p��ܬ�P4�y{ǩD	Z��;u���VAOٚ�Q��H�A#�DL�@�#�W�E�`����s�by���m(�@�v�k@� �n-J��`��4j\�+{�/�TCEǲ|���>Qm]�Ҷ4Nm�|1��M렏�G� ��?�Z��{47�1��}0ܨ�C�ZŃ!!Ӈp%U!'y���I5��K*�����*aė�2�3�Nդ�w$k�Z�u��'mB �	T��������GB���g���(4�����n�=:�bf��Em�� Q�Z��˷�������P�'�.H�l2�SgY),�H>�jL8 ?��j��~��u���b i�HCX(�R퍧ruPJ�#���h?�5�o���K�,����H�Cz�=�S=��|��	��}�i!}�K?���;W;��C�1�q))�(K����I��--z� ��a��󦎄�,r�(������Y����9ȡ1�Z�u�f��,��2J|@�+��2G��r��� `֖// o"60ĕJ����L��#A]�����+�$�c%���Q��Ų�Sq�cK�l����7N��3Lj�wwl5��ѕ�g{���Ć���Z��z��L���!�<U�/���|��wW�ء��CR�	R.7'{4�ʮ���_�@>�P�N2'(d# �z�Ľ�)�,����x�g׀I�:vg?��(���sU�h"zL�G���4j�>T�xw�WJ�/�ChPI����7"��,�Gn�ԇ�����}:d�KW�X���ܜ�j ؕ���%k�����jT��_�n����ā�m�@0<��m_�Fp��@�4�^�z��K�@����A�dH�̄�3]�eO}�3�ܰ�G#Dj��+_�����Q��Y]o�y�R���ye?4��>`mk����ɐ���g�T��t��S�4��=�'m3����~KyS����jZyhb�t���9�^4S�<����A�R���߂�sq��K�@@��Z������?�:��h�x����*��`���겞R���	�oǻ0ȉ�/��iz)sq��ER�MŜ?|��Ղ��輽g�*YԽ��m  �D.��(��[v[�,����9n>R��.1��!�Hf�&z�3�ZUn
� u�F�Cĕ9�ڋ�����XcOU݁�ٯSVh!������9J"��ٌ�Vv��p��Ǵ,��~���H�hRɈ���L��X=1�7��?�_|1+��,3�4gD����4�ˣ&+jh��[��R������a�o}L�Rڀ����I�kJ�`}�LV��>���Ѻ�OS�``�X� �q�I�P�]0M̼j�v����~O�����=�q�,A��C6҇�t�o(.[E��%2�&<������R��[,!�ώ�ߛ:ϧ�B���gUY]U������]o�AJz|1���4:$}"�9g�G� ���B�.?W~T� �/�Ù���W<8�c�}�|�~�J�&v~,&�ɕP�S�.fّ^q�̴F�fJw~��2�uo�9�D���d�m��{P��8�7x�Ĭ��k�UD��t�f��^g���I��'�ha��Y
7h|�*>�\P<
E����\���4�3%u/��%������c�*�= o �2s[!�W�F��x}�[;����� i��Ơ�Z�TO���Ӎ����>C- J����}JM/?��,��)i�?�>�%��^AL���+�pL"z'cbp���֢`�d[)�S���3�v��r�l���B�	P�"����ֲ��L�	oq��W��lw��Q��Ș]ZfN����A!�y�I��(�%������P�ڲ��J��Ț�������d�c���� ��@Bs���=ڕ�-b��_��~���<XX�e�O'@�5��%W����!��2J^��5��W89�l�8o ��6�Kj���<ڂ�4���q�ޯԽh"V�b��C��5���{á�����eu�3X�ˡ�Ѣ�i4��e��K��kj�Ec��`q<bM���ZKx�P��qN?�	.L[I`7T4lζYp�P�����I-�o�k0q���R8i�|笰-��N�2!��i]JbzgFK�����б�'7��D�֜��Sa�˱�� ����B@�r�	��2�}����nD��
U��5  ��t��<�j��ky)p��/g$������;u&���)SM*/D^����k�j���d"�/����^�@�
��5�ՠ��B(�p�|���T�ż��Ď�<�䱼��,�_{Ȭ��O5ϓmh7�k��N�\�|+|mo'������{�����:\�Z��F�Z��5�}�*V���_y�����yN�˩V��Z��,I������g�)܌��7����}��V�	���|`���MY����GA.�����d�������"���gBy�R�(�W� J��s���(�H*�mA�U��� �!7�Й�L�}ｙo��R��B�"��
~����!�
~�v�g>��x�<��V Cؚu!��{݅_}��Ճ�[K&����r��Ak��ɶ�;�YXN����4�7ow�ʛ��6�{�a��ů�<���P$�[f�h��;4K�J
8uЋ�]�,%���Gg��S�в���0������HX5��4���w ����-�����qk�{{��E�qo[S��8����pb����^,�jk᧖n�]�Ca�&˩.����ʊ��OR��k�!>$y�b�`�:PD�f�verg���0xPĖ%�y9��C��A��p<%��7�ziW�̗&��ck��g
������	Ur1���a�3*�f�ڶ��
}ʙlP��ñ�0[���,�V_��A(����k�M��^�*֑�0��:�E�Iο<���QJ�ƶ&@��`>v�w��o���=��w�$7�(�$��N�	p��L�1ޚ�f��`87e�V�a�Y�ei+6	��,����ׅMh��i���-IhsY�>�1�f4wF�u=�C���c���9��R]g`g���S�!�
ػ�H;���?G�fs�؟����"g,�p}�R��R�E�Zʐ�-��,�ci���
����@R�H�-�}�[9+�~=CȀ��(����
V�h�u��qB,�4n�����˝^��AO��Y��]o��C{�����4jt�^��L.%�j���}��H�Ґ#u�8~�Ì̷�[�g�~��M�2���} ��bp��}�;ߙ!gzd�����,�R��#������t��f+ÆL]�]R�@��pa��./�d�#(��{А���v�@�^�һ��5�i���+aET��H̖7���`� Z���Z�X^A{�g��{�}͐�BM��]׏��ʐ�D�,"-����m(&�rL�I1�,6��hSb?��*,K����-1��#��A-�����\�6B?Gx�6�U��_rt�v��s�L<���w���
3,Tr"�QG�ϡ㐎aǟ���J.).r�Ik��{��}Fݎ4j��{�]u޺ -k�rH@��!E��(H3[�٢�HE��oP7T��ʪ��SO��؃e+L�#~Qz�ud��M	?���ۖ-��u��a]I7P�I�n�~4z�+�Ͻ�O�5T7Se멮S�;�S]�Z�*���1�4�Z��`{z��� ���o�HmH���˼�S��m	g9���NWm�k���\�PP��p93hU�*t�R��k�ܖ��P� ��1��v��ϱ�BJ�:�攁=O9 ��F�ا�e���ǈ�fHz?�ر$�y���ɥ�DH̗Q{S�8>��;��RNJ/ ��-�ˬ��1=��h�u��GL]"`v ��͢6�k\�@V��.���d��OEmLB�Ҙ�Ȏׯ����}��l�#�D��=1�g�T�֚��eݤ�T�)��e�1��(���A�ZOʳ?o�N��C��6��u;@�~Sۘ!��ZT�O
n�T�� �"2%;��b�g�G��r8\��G]f~Sl��vg�i#y?���{�OC1T�@���c�EJ�U�u����@�]��H�_�;��_S ��|fŃB~Q��4F�۞��;��2����J<j ��3"�RJ��9��RK��d����c��=�\���@�8�zK3K}���̘6�-ku�+,Pi$6\���By�R`�����~��	���&dmP>ץ��&�8+E����[�Ǒ��T�4ܯf�*-�)|[F�O�jx^�~
K-(�ޔ:���G��6��7��bǤ�uJ����:��D��ؓD��k�IJ��,��2�G7��ӎ��/�I&��"B�jd5P �B~��a��%��t�q_�l��_�8��KCC�H5��E�'�k�{G >���q���Ġ���!��"Cp��~�T�F;M�����B�Ħ)�u�w/[Խ�1p6z����{F
���L8L�'&-~m�?
�����M���V��˚`�ٛ��X�_+�r�trVɲY���r.�K�T���WS=S0�r�]<�f`�
�o�|>��7cN�E���?'�Sʧ�SF6��a��4H�${�C�!!��K�vO�ݱOK������_I]Ӓ��MM�Aߴ1���"�7D{P���?�dHB���h�,��j��)��ܤ,XyP(�Z��>8mu��k��|=���Q@ ^�:�����7QM�Fb�B�c���'�zP��PM��E�8��^�V�"�׎�2�d��(�sr�-8�_�7f�
oS���;�u'C�X}���yA�,��f�/�n�,��H��	���!>�8�|�;3Ǻe��'�����3k��FXJ̩�r2�7k7���d�Mf	3�'�3�j:�tB��I�T��=���j&��|�d7���iW	��~���Gah�µcB&�~s�h:q���Y�~z|�w�=�Z1/l	�66�휮���v` �fI��ڂ8������f�NB��8awA���F��R�.:�!�n���5w��pzp���5�~��zh�(�t�H��T� Ե��|�5A��-W���F�*M�5/|���l{7���d��C�̡9k�}�]c�Y�8a�9����<��~�X\��&�j=���C�t?�"e,g>B�s���v�%W|��j�����ԫ~���F�=���?�.��7YU�D���_bV���M�F����ܔ�s�􇃑��պmyn��b�m/�� �\ӭ�X3�����O���1\o]�`�Ѧ�m�/@�6�����3��f6�������A���&gz�#�M6v��z���4�猟��߭��cB�y���X@�9��MΤh#vV_b`�-,�
�"��l��zUn#Nm"�~��F����������g�9�K�z-�^=�@�i��q�Fc�.���K�Z�xI��6Ku=��F`�g{�VD�fe��7�|���*<�!:�1�]�6t�}d��M�N���in�߈��Ǽ����&��)���w�3ޮ�Ps�j����'X����B�m\O��'i�>�*Jw7*C��Nvb�g�F���ו�fjĈ<�k�8�o'6� l�6*����\��9�6�'��|*腓�<���U	X�ٕ�N��7�C�+az+����v��a�+�va��!�a{��f߁ד�穓��=B<�Q�K/��MjI��T��|�5"\�d̞�)LQ>�C2B�$k�?$��¶__�S�d�#F���tɈ����!s.`�rvx��Ȉe�7$?.OH�Ųe��J�4��!x)�$�!�)��$��̹�Tk�!vYs�Ǎ���� j���Y�%�Ïz��h���4��2�u�괧,JbW��'l�lS�=�%�-��vϝ�aF)������t���1u�M,g�S�qLYk�R%�~j:u����v�d�Q�IXDV�����P�/(��M���燻!Ԑ�N"���3�C(�&(�>bV7C��kwy�ѨG��ȰC��l<�X��uz���n�����M1z�%��!U���\�+H���L�]}-�"ج���?%��Iw.Q�����K��,�y�e�fFy�wv>��0�Fs@q�#B��3��%G�i��Z����?��h��k�|���ٽ[{ɇ����8��⾵4C�����)>U(��iR�wA��	��:\�[Lό�j�:���a�xO��J���Z��l�B:�#�t���5r�ĩd_�
N�p�a�g��D5;��5�!!!���s�B�����I}Hl�طZ7�C,d����v�b�j��r��U��	ɻ�)���CaY3u��y�qz�D� ���"��w�����n�)�I��1K�]�e�t�W��Q���.4C��A���>ST�$@nJ_�Yf$ͯ��*,�j%�	���f�T��:�:"�B����=K���!9hP����� ��oM���T�E���CE��:q���\R>��{�&������JQH��H�2��u�DM���k��eWu� �Cbu�6/���
�nѭ��j	�[UD\�,�|�!�4�t��s���lT}��:6<�z{���/^e�# B����W�����~3u��?������:��AT���^��	JP�͊��-	������{e�C:�,pi+W�#�gh��҄,:�C�o��K�E�:�&L���4��10
�������Ѕm&ݞl_��^Sq#�c�0�b��u�>�&�#�O2����!��v#AjP_Ǩ��ԔF�_oq dP�,�����n��Q-�#=�6�E��K�OK����~��3}���y��(��Iq����`Ӥ�
/	� �Z\����'�� U�b��ߋ��~���nM$&�1'��P ���q�:��Ϊc��$;�a`0�_�5A|"��?[=�6�}g���m[���E��u���4�8�;���@5��?U�"47����Y��)x'�iBv#*�I(g� �<�����4a�`j������ �e�I�}�_�o@LY��w�?=I��������VtJ9�j����(�ʓA�<=� ����G�%�A��;��?<f�!l�x.�o�6�u�{� ���o�:��UgZ�B*_H�/Փ+NX������f���� �F)d� ��q.����F_��Ҏ��R����aaH
�N	�]�
F�l�~�-6J����U����K�=+����"�E�&ߚ���ʬ��謬 ��G�,�����F�P���5��I�o�K~�9��7�G��)�ᣲtCm�Ҳ�v<h ����v��[%����M+�`'���%BG$���R�Z�b݆9�w��p`������c��2yLie���l������΅g�:��Ȍ�'\� ,|"�J�3�0��o�����-�*�б;`&�t��h�W�ţ�J	!�(&p��1�Ы�=�ԯ���ϵն��2���L��ݧ2�G��L�ѕo�M����������^	Q�&�袍�WTڨ��w]R�H���U���-2������Q6����V>f�q���+���g��rf%��qew�I��,����B	�)HY�K�1x�b�Yڕ���5�W㘹�r]�@r�}˽)�J���@@����JL.8B߰�li6����EKk���N�8]	b9F>���V)��]��}t�\�>�E�o𵋍��?�{� b���p����CGJe�⛤�ra�bw��Z�t�Շ�7�r��	���}.Ӛ(�)�;>��bi_��0ɘ�@W4ݨ}/.�Pt��f�O�k�����E����o���r76�M<�*��ꟼ�<�]��̊B����@g��;q~�k]U`i�$�o�P�q�E�x�}Ġ#tt��dm�i_�9V��r�`2��*M�Z����)k&��a��[ܤ��4t �� 4��:�9������
��M��O�@\����3��b��Eb��Q�k�3��82T0���*/��an��/�PwtZk��^��g�C����%M��N:R �e����I�oҦ|�E	Sw��cҝS�.}:�௖3@4����^��4 j��/�:ÿ~���W2R�~x�'���'����� P��A��N�U��
�{+�!�P��tۼ�ך�ť
�[K��y,�h��ß꒎FYC����P��D|�7�?���	���,z��t�u�1�Ӵ� ���a e��
��X.T$Y������Lط��b�r�6��#��4 �/��}�����;�R���?(9�A�kN�?��_���ۅ�6�L���br�!.�r�����H�-����9T�W����/JP�g���ܔ3�a�M
���M�6;��(�J� �	�r�5}��м��y����E/�z����I NS�%h�J�,hY��" ˗�����{�3�[L��QCY��alhJ����:��Φ5�b����J��D�-E����*a,����K�bnK`$$F!�X�*b���������]�ZKr=�n�(�,��[Z_=b���7>qL7�,�6�X£���^F&����;�H[�4l`�ΓMo^K|z0l ����K�5Qbph��a��]�e�q���ۻy��X�(�[�Lk��FQ�J�