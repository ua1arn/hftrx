��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga��ʊ�tl	]�1�f��"�~�őᨘ��+��-��&3rLTf��j�ս� ^�]�)f�.F�_u��v�7�ن7N��[��j�d��j
æ��v�G����]�&�AW�2�΍1��B{�G2����Qr0�izC��p��%��.qÇ�ye2Ǽ`t��FpuV����A�\��i�I#B:
�8f��
�#�y������{Į��S�E���Ų��:�+�<�o�����*��� �V��a��Io�8VHHf�1�0|�[8�f"�-Y�w�
dc<<�K�&��o��Ɓ{i>��P+E*����~y�L��a��|�'5�qe�U���b��tmF�m�����M�n�6G���@z',��b���-���D茸/�
b���!�*�������I�N ��.�J��o�871�.!:�R�
���r*Q�����c�~�T�h���$�^�[���h�_#O�~A����΁E�=\��Z�국#�[AX�?�ρO0���������S��Ɯ����\�"
����|}��#���wv}��S�tW��l�2lN�=�̈򨕷��ZR
n�����Gh��[d;��"�W��c��K��'{���+;y�}Z�t%�؉��MOL)�[����'�U(��s4P.3v�s]u�K�[��_j��k.YU�=���R`E��H�v�i����Z����!N���F�����/�:O4\Y��wP�}���7x��-�O��6t��1RY��w��zU���׼p�6qj�酉)�P�U�eꥐ������}Yx�6�� $����GT ��0�adK�|��A"��F�&}����Fwr��uQQ��p���;ڗmi-k���TQ�	 T�&<b}���ͅ�n!���1�{�cX��P��5�)�H��ggƟ��PK`�����&t��K�de4����qqtvuI<�I�B^`� �BK+��;�G�]���xI9~���9����Kg����7L����ߐ�4�)8�w�I~#�l'姅M�4f�e��K���?�5+��j����&�'Y���6g����������<ݮi�Z�ے���J�\����V���+I+@�\���c<¶�<�5���2�� <��s�$���]���Z5?�*d�@�l��gC��f7}�M���0C�H�D�Cu�S��G�\~y�*F�Em�M�ҹow��%��27��	J��� �~����	��f:gc�
{�������U2��X�꼟�<a0=n�Z��z��7E�9���]6Ec�=z���~�'U.�:�I� W^*LF��%k)ҟ�/�g�����Z)h2|
������2k�ۯ���{`)#z������T�Q �l���.O�;4 �\c�Ui�d�2���)֋�ݲJ�G������DP\����&�4�'*�'�jy-��^ҮZ(qC�PRW�;��ӛ���($�̟�_��5R x�|âpX�Z�}�+�|1�q�d0�����Z�h`���``����E�[}mr���~N�����ty��ׂ�a�o����,�1�:˻Őr_�
%K����l	��'-k�d��HJt����y6�?��,�.ኴp:�H�]'m%y1��R�r7M@����q��-����S���YEJ|�ݾ�ϲ*~�u�*��.)�GL�����D�2x����ˀ}�UM�u�Ė-�x�+�皞�&���7�Uiٔ��Ў�x��SJ�L��w�6�^C�:��CmD���L´�DtW#�N(K6�ޡϙ��6��d=��硉�W1�Lן~�r�~�;�)h�pM� ��>qX�b���ψ���|���u?M��8�	Z�J����*}�D��*,�z�Ȓ�W18�����-0���'�A9	0ܓ����!;#�̯Jj)�L#���Ԓ �y�����}�Ìo�S�K%!�>@��<:��Q����(��E�`��B�z=�aU�W��>ߺ;�]�,,���o;�P�/�� T��<V�VrH�C�8G�ȕ���y��`b����D���������8��z��1�K�S,v]}-��̕6�S-~.15W�<��l�����s5�Yt�ץq�����0�p=p��K^Pa�����L&�f�a^������j0�M����)�z;�f0$T��H��٤M܏�3��%�a<m�^��u�MW���L'w;@��` �(�B��L#>fPAI��@,>�Ƿ}�%�d��bІbO��ax|):��wu^m�!�������!C#^����}��c�<�s�KNE��ءg��I�[�t]D��$���%������ݵ�D&��@Pv�2`�j�Q�e>�j�\�ygB��!x���qZ���	�~�o�Y�B�oͳ켾!����`s�#��ԡ�L�S*T�q�$��d�b?qsi}��7*
��n�� �qCe$̈c����J]��q��&	�o�EϞ��g��)��%�FK�=v�U��{�n%%&�Z�^�`^�M�i����'?,`9)a.:�R��	bP�N��x��2b�a��r1ŏV�H�>�^w�*`��c�d�A�CF�����q�d�<He�pMiCK���|H��!Rd�I��Uf1>�/�'n��a�W�p�vܵ�xo!�yX�X]H�}U�x4�o�������a�!�K�\l��G�_c��)34��H#/��]I��6�3������*fH���e,�b�wl6�� �Wi�c  �L=�YBO��M;�������e�Ъ�5�������u�JS4��T�]u��><k�	�%�i!�	]W�.֜Iv��oJ�{^�%�+vo�YI��֟5\k�{��]�`���oN!�sH0h,�uꓟQB6+ioe{E3+&a�d�)�,R˗oF{��ν<��R8�K�ʼi��L�9&s�I5VW�����֜S�}�(^I�+G����Ƒ�6�1Rz!��k��Z�c���'���&8��1���n�|�Hl0q]�ٴ��9�������_^�s1�����z�e*s,h+�@`�w=��������8Hw�����}5��	2/I0�p�9n�	}1+<�2�ט��K������3[�����'k7�N��W���Vo�g2 ��9-��o2[�����
��w���K1]��g��k\�D���s&�X���oaO.�"]����X%H@����1T8�aI�!v<Μ���C��J�Z ���1�J:X_���h!no��$�u��X�7��m�ؔ��A�Ö�[�ڈ�U�O�@���AThU�����ܶj%�H�3\�8�v9�!���p*�b�$�KC���[�1����.nMb6�%Lr��g���w*	�>���R�q�s��i$B�-Ҁ&|���3_��H���B�`�̴����'*��eORJ�A�AVa�aE��/��&�H$���	b8��.G�rܻq�iL$Gw��aO xj�/ ��1i��s8����׵��؃�GZC�L!!u��!ޯ2��h��5�:��D|�y'�� �����5��À�x����p%RՇ���
�n����Z`@Kw߂w��.,辙��^^�l�YFՙ��0�K]&\ˤ�k�J�g�G�����#��؉���M��7���>X�ȝ����5��fm���L�@ٙ;K�x�j���3Cr��8�f��Q��~��,8L�):PH~+�;L�VK-֣�x	�rߖ���J�(!aB�B��y�������M�#g�e���j_d����#�l�ȔSŨ:��ᑍ�!�����+('z����l�+>����uG�T��X�\w7r�o�}(��v�]j0�4�K�s�����ee����T�9�E�k3��ۂy.���NpK)6�&w�<t;�$��3������V�.{ws����G���3���<C|�6�[^蚝dL�XR�B�1���t�V%�̊��N�#�0yǂm�+�4��@J�=�op�G�r�P�矖&
i�\�`wD7~���06��Ό	=��}UEn���Y�k��@Ü���>�arB�\�
qC�-���8P��(DrE��!!�ĉ��q%�.(�%X鮭�����~�mXI�F���Q6��л5�&Jĕ--d�(�
�r���@ET�^G�7p���u71��۞O�I�A���M����/1)�������F-mԝ�������֨��?0ˡȍ&�5��m���eJC�s��2��}�]\|�E�bb"���Һ�,��Έd�D`����Rb�h���g��P=H&�ׂl�4usX���������#3���@�`�c�*�8L�0k1��q$k��jP�xǅ��9n�ah�{*�Oyh�B.o=�+&n��N�s���b�.��$�5����z� ��+gFi6��]^���6|<��.9����%=��D���D"��Yd@:�*��k�w�I�B}�'4kx�#���[՟ �J:*�>ϭ��F��*�x�/(���[�J:d46ep/�3f��uH�S+��Dv����=��WZ[~|jG�Q�̾�)�}S=���Y�\]�\@����e�f�/�В��J+�	���ү�Y�\�P���)N�)���[f?g�g���I+���C��g�fWZ�Yn��а���iSp$��f�` o��7�p��ч�L ��<.+^��gI����-�́��D��PAԭ`!�u<&%9E7�����y�fŲh󍫥̈�,��E�X��r6/M� �OO|��xz��-h���e��pISb�7�,�|�dJ����:�p���G"��[�������[��i��JZ�|�5\,sQR��UegFK����8~
7l�4�B�c�cs��_����ܞo�(qYm�\�{y��:,���H�(>��d�ؤg�d�/J��>�>2&5zK,Z@���?�	��b�\��h���#��1�8��}kh4eAQ���+(67h�*��F�|�O�����D}1���W����)^�@���Ie�?����m��H�z���P��հu��͐�dƀ��5��*�Cb�H�g[����Q6V(�)SVъM��?��̜��&{�.�jf8[eR���r�%�3mjz���$�X�!w���I�+������<�U2w\6;�2�'=�J F�����-�W.�z��;	/�� p����c�<n-Di2h�<�{��7n��+�z�S�n�o��K;�H_��]��[�C��b�x�����MA��QMG%jFK\� ��{���d
(�Ćͭ�X���"ܒ��늛�T~}ؿ��q��ȗ&�V�0����3S��)�T$e|�ʼ� �wg��dh7��  �CVmt�e�3}G�*�K���<�7S��s��A�X��z�6Z��&��x�4x�ml�6�NSb5R)MAI��"����X�5�-[�M_5���,���Lr����?��'�M���zB��׈ ly�}�S�����m�_��]u$ƞ��
��'�X�A�5ѣn��e�x����R��;g���R�P�2��#8!$�y�SAb��IsUv�@W���ZZ;�=q��ʛ��^}�a��%[?�/��ĉY�;�oj��8c+���+�r�d�ǝ|���G̍
�h���=gkK���~��N��J��Y`]E�8��@�	��덝є�=�]t���s�I���rW�o[�� ��Ӂص����-�G�;s�G\�`�����2E��(�4/+}X�ӛ�O~2��/���W��Ewjv��i?cL�~��s�U9i�?�o�ӆQ���5�[�f�~��^�Z�Hy����.���H�}e����9/$�`��4��L�Dpce����ف�����ل��Y�oz-��Asm<94�fd�/[�X��Xx���P#Oۮ�n�	�r��8��e���:������_�i��̩����<�.�`ҭ�O��NQB�����#��Щ���!����S��EK*�4�n���½�7��na.����y�?�=Z��jW�d�^�sO������8[��8+�}|U�G� 5��IZP҅�(��j�Мn��赤U(ZÑ*�iR�ʑ4\E�	�4����<V�`�M"Y��"O0�uT&H�~���䁬'R�Р�<L���]�(���ڄ~B�J+��I�O��V�Gn)�E]��@p_s{y����� ;� ��_�s��d83��p�+�f/w�!;S��C�Y;A{���:v�M�֜���&�$�o���[�© ��L$��찪�'�J�M����e^�� -'�Φ�x�2m���&C@Q)빥�yS�DNul�q`ϺdK{�Y<�b.
F��[���^�#����![�Mf
)��shHM�TV��րֈS�b������l�w�{ ���w���$�`��{eW=���b�,$�A��?�� %��+�?���GHL�ӴO�Β%�͉N	y���&���#��
^�J�P:"ؘ����ׁ�M)��LU鰤�z �9�2l���i��`�\o\� N��M0�L��
�w�Z�+�W&�^������5��VA��E�&h���;nS�.�խ��E���#1��=�:J��WM8�^���;�Ϗ�[�m 74�q�E�G>�[w>���������ڠ��.��?}���.Re�mc�=�~[A��O%cDD��<��V�J"Z�����ϛ���L1r\�y��&s���%� jj�1�v1�, �V�<a���O���e$O�D��	�X|�K��D��(;�H�zM�b���(���8w�{2���<aA��ރ+��$P+a1o�� 	���v��YX�/���T��0o(,	��'��1�.J�ȿ�z���H^s��]mc�M=��9�r�b.���6��.ˍ}tP=e}y~X�O>.��[j7n�ա�rE����̤Ż+28k�n��	�g�	z����L��b�4���X�Ƹ���i�fBWi�ǌ&���O2S�����U@'���N�S\[Ź@nMI��I�t����&D��ᢵ�jʜH4�E��R�3�1��s��ƾ��q�`�W����=9�;��d�]�lL��6���6 ]�I����ȷ��`���I"�i���U��d�UOpع��0�f.�dR$��9�P�� �ߛ��kY���/(��;&ڷ�8��qw�����V������ )������-�(i�]��,r�I��P��QTh��O݀�W�J���l2����70C@� �Q}.�MC^"(Z_ l�ė��T{��VM�^� z!,A&�Ti����'
,��"W��s���剈U�h-���0R�����0),?�D6�<<}�[3nB�	�o�T�z�!J���
)�}�������~G1���u�,Kp����*�����iP�c:�8Gk�q�I�^8
�8��x���i�R!�b)�ۣ�qg\�cZtW�5Y|���Ah���?(y[p�������.�ѭJ�T�?�_%�C�����V~��;ϋ����Ј��R�Ϯц�)	��M���\�1��<����R-�^w��4�R�6��gz��}������@���u�x �c����o`{x֚�[h�Y�w;�r�"8D_�(������sw YL@?�QB`��n��"AG�JKN�e���X
2K�+�Qp�݃&�I/e4�W\�GG��������qw%�4��`	���L�yqJ+|l~�v���� .D	pb��t;ք3��:�r�%k�n�Y��m�+�`����Gj�+�7I�[��w'o=�3k������E��
&Sr+i6��O���oN{0,Qt�D�9I�L$H9
���-����]����?<��}oi�HF�π� �_��;�sg��b��7`��B�������[d��^\�5
��%-��JP|X�m-�ˤppς���{��*TS����'�`9��������|Lb��*)Ѡ�A�)>��7l�&�5��@K���;��aR����p�]��Y)�V��h'��Au��r���&ʓ�[ �1*�k^�1�"�J�>�����8��E�/�K��=>Z�_1�R��&¢�ɤ_L�x�Nt�$f�-k��� �����tVdb#ȳ�x�@�AG�� �!>.�C����+$�|��׺�mނ�:�i����N$�#�ǿ�:���'��
�P���A��,��(_�	�������E��6���<���G��'(��7X�Fާ��Wk�^1��9"[Ѱ��w@��񆇞�7]��X9��+�46q��Ђ�ۖ�.�O���;� �T!%�믙���C�y��qṬ�����;:N�	�8��:z���xĹ�I!��&�C��z�M]��]����*�0�d��@���M�~�F�U�A��T�j�\��c9�V�:ϸW�~@x�����q=o���W��7t)����}���sIm�'�X�s�����N��6A��͵1N�QE�uH]Y�!E���5r�)��7S�PtM1������,=G���O^O�蚑!�nvraD�M�V��-��i���j����ލ���p+�tZ�A�G5jR��VÊ� d������+}���mъӨ&��}3D��{l9b��.�l�ř�H�e�*&�����5!�_�f�����J�蹡�',�Ye���ئe�QI'�_|@Ǟ^��g7�~B��(���|,�L*Ws�C�rd�:����ya3�q�
u���o5Òg�\��%�h�1Q��o�kS�|]�.�,%@E���b-��R���v�����m��2 L������I�vb��Wu�Q:T�L����C��ZXY�E�}O�E����*$�9��M9�'����^\r�o��SQ�̀!:qAsڿ�PN�z������iҋC�ÃGj��HH��5���E#$	g��Kʩ]�DD�Z-d���wW�8�i!w��w�7�d�J[^|���F�)*�S�0:"�'��O,wƪ�4x���Z�(�C�S���PӒ��t�g?s�f)֫�Q�Z��w��9��h�� &f? �m��4C�����V���d�?�̯A���Ğ&㡔NRmv��vm��4*QO	F�3�m�ȑ�y{ �9\)��(i{*���Ǔ?y�v����q,ft!�Io"G�u�"�$h�$��d2ڿ��_�	�v�[k� �K]�>�8�7ߏ�EZad�����k��$V����Xs�G�_y����(�Uꇯr�z��F�H��n�N�	!z���7�����ɘN1�`:Mv#j�S��Ȑ��1��|����+�� 	�k��B�#���'EGB�t�����U~�y�����{���%�*+�1�	��E8�����`���C"|�Q��t�<)�l0��SX/���lj���NǦ�T�Z���$�Գ��+Pw@��ڣ����i��ݫ�7]��v5���U�w|�$Oi����@1/"�{#(A����W�(���Tc����`�bՑ��JC���ݕ���mr�x[	ӸC�x��m#(#�<��F%�3(�cc��$r�Gۍ��'7B�$�+N��bf�+䋋d<$�DA�!�a� �f�F�/���KoKm�}�U� �ˊ�F�Ц�v�E@ZOL���D1>|\d��a��f}J�F��� e�!Ff¿�����h?Tq�mГ�&ao�"�ѐ�Y�\Q�31T�������BEDΒJ��4�%#È���bY>'1\�u�Aky+,���om�`����Ǜ��tjބYm7G$wʀ֯x��qd+�ɟ�7U�ii�3���~R��:��s�h����{c--r)���,qTv7�3�E%C˼UV⿾`j;�r�]>�om.�z��B�k.�H�9��lkƕ�y��V���4��,Vj��1bެ�Ypج��_^9N�jjrm{4U4`�2�ŪZJ��#j-1�o=hq���n/����5��:}1Pxq��B�wJ�m�a�c^����y�l.��>.�J��e��O��=��,_[F������4Ϥk��
�32��c��]�i���H_�5�q+�٣I��d��Sc��=2]��/kqS�7	U38���w۱��C�{z��}��R(��ƶ�ޣ^�J����^����a$UMʊ���ц1G�]>��˘�ثwT�t3�I"��SD������ٶM��ƾ��#2$E9�'0zK�>��&w��ڹ�k����X<PH$O�Z�������^i0�Z�Ѵٗ��ⱹ*����W���j�Vk�����۳	0g؆�S�f�KkF��<}a��c�>ı=h��g����]ޖD� S�Q��?����)	 }�}����i��s���P�{N#$�X�>�$���h����Jޜ����g�i^��������Y8�3W��j��:2�zVeK�;�q�C���p���M�p>:����.Sa��1"�zF�� t֫�|�`陁������ ��F���P�(��HhG:z�s�MG�x�/K�%�o�Z@�w��$ߐ� Ovj�a|f��arc}�Z��ӌ���5�0��}q���/t+Jȓ-�=�����Esw}��#�@
�AJ�:,;S�z�
l���e�^�*��g|j.�T����Ԙ�E��?Eg��4,���\�SK�hH-���d�s�ulh�#n�4M˧�[탱KE� �t��h����_��A0."����8P�\���o�=h�p-b�����.� G����c
(�?�A���Ԉ�̗0{�s�ٙ�4�^jotKu�^K�}'�g�ܵ�tt�7��1R�玨Z�[L��0��)���mX�\�x�r��ȔS����>	.cs���E�č^��lD���e�м�����~QށG�V�&-�	�4����l�2S�����Yy���L��>�/R�owЀ"!�z��1>�VJ����-�����2��%.���-��z1�@��)��HSd��jY������D����M	f�L�c�{B�"_�3$�8����Nؐ�Z٘��&5�̼T2���g0f�U��@��o\�"l?�x��چ��~�B��zxxGfm�ja� *�uYr?���р��_�n6n:�������/O���3��ԝ�H���&E$D�!�,�~�ʉÀL���΍�`_,�;_W��-F�l�R,�$l����epNN�^�.�6�l?`L%`��ד�6��k�]ܰM��k�ͭ�����bg̏��s�}����j�_���rV�y9��	xD#ۯ�IޯU��x`7:� ��r�O�=,��~R�˨7�t�M-b��@Xw�G�8CF�ת�?�<�%�$0����)�A� ��{�~����Q�p�1�S�Ǣ���w5{..�Y�o��?d���*-)�\!�f����}��j��]�(0?��Xq�t��|z֊9��bZU<��B��D�[ W�x��C�.n��f�A8��ݣ�=�~��W�ߣ�J������X��WD�I&A� �H	X�bϿ�H�y��cG ��N{:�ZD�ꖩ����o}�'��;�[�?Y��/��>����Z]zk���j���Dl���~�n��'z�~pUu}��R��t
g
���n��>�O������^�`��U�x��3"��}��)��u��0[kJ�\��bv9�-h��`
��L���a�G�F�O���� <t'���������� o�㣠����Jn��,-��N�y>�a�6���g����Ԇ ��*{��/��:&��6K�^�r��ˡ-J����Pu�#�m��g)Q�s揘�A�:̮�B�t(����RM�`)hNe������e��P�i���k��Y5��G�X쎭ǢrW��֝~��}��.��i�ڑ%ij�r�wN8"�̞Cpw_m�v���
XV; ��κ0��Kگ�x��y�^��2�<�H;�U�_UY�Q�T�?�E!�
U�=�4m!������<V��gr |mc�G��lD�	�+ՠc~��XS]�_c��噀���7آ5�L@���u��:(X8Y���OM钲�@s���=:lpU_�_�}Z)���b���&ohH�`�rI�G-ϠR�S')+�^�}|]�5�.�ζ�9>�����	���렩�b{Q�Q� H��0��qa0�L����n�K��ub:F�d�4��F����U�"D��V�t�(����7?�b3k��(S��w�z>�9OlV&o��#l|���6"��xF�6�
�5q�x��}�bU��W�t��qA(S�]�8;�:�Sɾ�m �;c��Q�
H�˿wdS]�4JmgFU�]�e�Ac���?�N�
K��z&�|P7��&����+�G��"$��?�����bem]�Z���������H�CSr���_��X�m.��u���M�<4��-b�#��Zb}��	Ղ�	`/����o���Im����#�G����K���8���/Q��Rn�
�bbīB�K��]��!��y2��<ay��=�����m���r�Y��=���l�<'x��H-�.��芁�����8#;4�]z�l����J;�����_8�8�,����S��
�R��"9c�ɊM*�?eth�ᛚ��2N�1iu�h�����77Q����q��u�	��ۃ�JI�!�߆��w�2R���l!�j����_��2^�3���$� �}5�"���L�-&�k�Y�WZg.v-r&�+O����\#���`l��`�9���-��┬ 0�պ3f-M���:���gu�:�,I�ϟ���;Ǌ��4���* EI���6oFn���3���eh���Լ��X|V�_�������;�HE�)&Ώ���0-&g��b9`�ͨ�����֍������UN��;Q�����B3Q�X��)��:m��2��*^%0�QĘF�᱘���Ԅ�>��^��
FW��3�vk���_��x�}����?$��ݾ���>r��N\�1o^>�T��{?��=�i=�Q�n��s�s�tLt��.&8`���W�Ȥ�#Uyo�C���5a�#I}��� �EG�${z}G���� �j�pFC��=�	bA06(ˍ�$���[���p~��Z�@遹:e�>fM��dq[0��i,��{�vpA��O`��,č-��y�HY�83�s;����w��ogH����P�|����3�*��%,�?W4:'��=�b�Z���uJ`n)��R�r�N�M����IЙډ���4�m�E��U����<;���P��Ⱥ�
'���/&�C���Y|X�:^?t���ji���XP�(�Ç]��̴�`�����̌N���M�����#�u���Ȣ���Ǭ�'e;Q�%������ƯB��un--��Sg$;E\����Qw�ܺq�;�,�wM�Jq�K��w_�����K���´Mޟ�|����Ӓ��jh�����<S*�����^�NQ>	�.��\��S�EF�f]T�Y��hn~r�¶���^�ZV?o��`�YީeE����ɼ�c��P���p|\'xջ��-w�~�ʨIr]fd��D���{{��v�}�d|KW�(��\�����]�dR4�ܡ}��tG��if�>�� �N  	x�"a�e�
#8Hk(�{�a��ȯLD�2��1t=F��l����*�T�])����\NhE9E�����b����z�(i�տ����>dn�N>�q��qA��lĶv��ڈ����mƓ�] �b~l;��5�tUV�g�����-g��F!���A���{��"nZ�)kN��@V���q�n����3o}�m�� �I�Q
���w^/6/�q�@	<B�]5Jt�LQ�ڋ=� �D�&4�&ȸ� �=/�}�ܥSJI�Kt����}+MY�,=Q�zu�����+�O����X�-t����W'�a?6}�J>��&��ؼ���n�i���Cwq܀���0Ci�����x��khC�"���4I�_t����L����c���	�(���V4-(RZD�ku2t���Ir�v ���,�Kd5�
n���[%$�?��t%"5W��Llk?��?K���2M�Ͳ�K�JٌPix��J�� `�%�z����bSD	#5k�1��Ior
�_�SI:v}���Hy�rb�""}1L31t��d��@�l��3�Q�0Z��JIl=j������{f�<m	%n-y��<�1�4��\ytE�ח��fPA��&��0z��`�d�@�KLuY�
N%�TBi� pC?I�����;e��7�sD����؞y��,)�z�gOCR���@�,�!�N&����+=��J����T���vL2h䉤��0��|����m���(�(�(�AΘ(qZ���2�?
�J�i�i�@���6�ʫ��tk�m��E$���ۈa��#G��	n�f�p���B:]���dǒ�h�j;��GIm�������?	�Sl'X@� @�#��Kx�;~���Ks"7���"�AO�{^��~*��.��On# �x)(R걯�oԺ�>Ρ�¨	�Š���4�gk����z-ދC
�A�=u�enwˉ�W����Z��K!�5�6(�E�4=��0ߋ�a�ч�u^qa.��{t��W�Z�	�ȕB���A�/��`ٔӏ���GحX�;���rLf���S)$���"�P��0���JJ�D��w��P��ZuhP��	f���dc'/QUB	�JjZ5�)X%?97����%*�ȦI?����^��5T�J�U�V�����$�������C9ms,L�/�ّaC��ް������F�q�����_��? hd���K�v���~�-K�4/~Jc�l�GXP깎���'��A^����.�K�$��*ӿ�Q��%x��x�2"R��S�{�zK�o��|ʘ�v;��o���9�b@�B��X�y�XZ�ROt�N�����!m�<��K��Y�%<�^����#5��%���ر8f�S�{�ޝ����io6�=n�>g�`ո}���� z�;��ыC7Tu� ����!r(�������+�A�$G7���ya!o�)�ٮ�j�V�]F`s��<5L�`�`
4�5S����Ѥ-{�\2��G4ҝ0��e;,�CFRbn��2�NE@J�_o	G,o�A �o���S����1^���@w-�q4�Hd�����k8�52����I� ��|�.26�pS:��`lx̶�k�uFTa�C� ��'R��3E%�?�،O�`��²x)/_G��M_,~c�Ш5�^�����Ի!@9��.Y�/7�|��H��t_��u���W���	�'��!e�LC��ź�nx5�-�LF�\P�m�/���	��My:!���O����4��]K7i]��yv×hg�j�K���k��V}���#q6ńQ�H�.�Y ����DƓ���q،Xi0�.�������^�a�`�]�٬�]�{ �c��S��`ۥ���n摷�hR&��g\Im���{�¶�
�`�u\��q�W���ĝ���a���=�6b������ς���<UQ��~�q�X�rp]��_���[�B��ðd����rU~t�s�)��|3G���+��h��P�x�F�>�H
�7�Lw��Ev"UHS7�M����ҢZ�1l
R���.�	KS�T�����4
zK�� ��Ϗ�,$����#��D&^��[�s�M�,���� I����&MjI��\��,��A.b�i&\l�������sԎ�rd��ǵ8$bѭ�-�]��{ʆ�����cD-(�)�����4`�Q��5�=���J�q���ܯ���0�ޱ��y�Q�x�>�)��r�l�Wޤ��ԇnw��@;���j 
�O����(Ȣ�_�*��ܭ�o�;�
z����=�����6���P�@
�؎�A,�Wd�qh�;'�3�>�o�uDoz�}c�|��tD�M8��d�{|�`�|F�%�<s��Xn�"�a: ��}Q�*��P�D�=����)x�������T�Bu��Qw�g_)��4��-��p�6w�I���v0�T~\y[���$����x�z\������0�#���^��d�L'�S����Q�v55�F���^%m ���}��h�,�����1��o��8=�Z𺘆��JK�'���T��B�/�Q��+d|���������"X�p�7���:�Q�][�D�M��5���N�-�a(�
+�Cҿy��������J�>#YY��v00딅���}�m.`rY|SA���qq���p�臡s�pӔ��c�C����ӒB&�k���μV�Ϭx˱�'�'P��N�lː_c4w����A�O��j��z����&b��K�zn����'���(��>̪ƈG�X�n���H@]����dt�)�`�B:����}��5�_����O�{����ʯ����T ����C��T���u�$��>�US�[�Ie�'D�!6�Q)���8�\�)>��a�?�쎛���ľ�ɨ��'C�*?p���&с���Zr0�`�֓Ì0!�V��W�bk���BHY.K i��1���%x�v}}�E�W5׃>vx�&Q�����R��.I�*-GI�-��yz5iy|�o�.�8���C�Ē�SBS���Kɡ0�%��.X��l���Bw��W��VGv9V�M=*�jh�B�:��\�>���L��L-QO����u�Kۅ^�^���a-ʸ�8�c9����v�[�|1bӎ�|�H8O��m
L12Ϭ���U��*o$.%T����V4�6��Z�{�����7l|����M���0���_�/x�@15N�!4��<�qP��uQ*�쫻L�ӿag�q��?�����`*�;ی=�7��	��u�9
R��,B=�x�d� ��&��	4�m�S=9���E/;7XUg�� �0���`����$�d����*Y���R����������X�e�r�+�4����Ǻ��6{054�ɨc6u5cX�4�8$H�F��<0#�p6P��$P0*Ȥi�M�*��ﶺ�K��w#�� �{b�"�sCDH��eh��-�V��9I"�B����d�H3Ìm3�[&%�=�H
���cp�Ϋ��R�T�����͞0vs��J	��x�L2@��#�JD`�P��!�~�D��Q3C�F\�BGM���M^ţ2������
3�7�쥑~f��s��,��O��~!��x�n��1��Zx*�����xǅ@��G�$3{�Pp.�G�.�D,K��ӵ�B�W�[���2G\�z�b�&�2��~�ꏿ-BYa�kU�r?��>#,�(�w�N5�$Ǖq �/���Ҹ;h�t�Lr%>yl$ƈ� �]x����"�Ԕ��u�4y�����֙��u5(Z�O:� y��t�dqW�?��1��T�2j�M����&#��hMA� ��P!Mq�-�Cj��NeU�ō��$s��5~����"��3����l�S��8i�N-Kk��K�JAg2���r{��׏5��NP#0,'qh֦#_f��21w�o����=
���ĳ,5j<nfQ�#�X[��/�Y����E"R��/�oѶ?m^$��m��ȫ5Z�j.I}�as�8/����S2Y�s*��s�
� 	���?�I���.t�{ٱ���'g���LʵC���6�fe��<ӈ��a����}p�TdN��cTr�b��)[�iY8�Z��m(�0�4K��F0�QE�ke3KI�aƍx4s9�̛��lj���b������Ea*'�*�g-|Qy~�����ą�?�ٟiR�0�U|'g5��S���wK#sΦZ�)���j�o�DsI�Bф�-��HGUuޱ��7������(j�oQ#�ȳ3hvNBA�y�
���xM9l@f�c+�j�<>?Q�;�c���h�����If���+�#dafQ,�@��;��;�Eh��L���Ŝ	�}����%2�M���/�%5rYz!��YC�K�@�&[7��Q�D���Z�����y�������� j�𣛌>GC�l�y[b���Ke��%]��w��bwc��m��������<^~�DU��'WE�N�W��D����4���A�8�V1$-�y�`����˛�|�6�h�f%z):��pzVvA�4*{>�����Z�������ӳk1e�3UR���=2�(�wPn�G�ɰ.*-ٖ��!�!�Dy���'��%�-����w���ߣ���'+��
��i0���|�'�t )�Mw�!.ŝ�� ���ua�+QPL�u_������b䖔��Z_ `�Ak*DZ�l���Z�{��jn�=�!:���N�Q�J%�V�T��Ć���b9����p�����_�|$?���b6��m��D�3@h��u@[��]�dH���d��͋�*_7;A��'旛4/��\��4!�UW���"U"� �4�U�2����Ug~sS��ͦ�Ck�m������M���~��� �[�~'^�MA��Q}�ߞv��Cr.��}&F�N��ֿ�P�U1D?<��@�w�hY���Z�� Q0%���ŉ;����C�Oߛ�/I���A��"�cv,�[�+0g�2�&��ICΓk'^ll��)� �/S�}Qu��]�%��Φ��B�0Ǧ�R�r�G�8f�~�{��'ڝ���)|��|��D��$���nθ,:���:�������9s�^qrW���dY����Ȝ���}�M
�%/D �N=X[�?L��	��d��1���=7�$�!�X�	����z]�s�D�
'o�ḣ�P%n�M�F�:��(�_��l?�߃��r�ц��k#[6��է1��j���CR$.ԕ���%��ɠ>B�l9���)Ǚ4s`�F>l�UG�D�࿶�^c�]y템�p�눒Ѿ�u�}կ��v�d<��- Z���/k��8D�˛'��EC�[�?�ʾ�Ԕ��!8r�h$#Fl� U����#nB�NkMv;�͡�#;��B� �+~�-�☺�?�o)���o������T#+�Z`�x��,{��O핸ݙh)Թ0�g�/L�>*��/�ר�"�D(r�C���� Yj�?ى)#f��Pp��zk,��Y_��Lj遹\\�B��}V��Lv��6���j����/+�����*�g�l�p1�j�:�R�H���Hݿ�R�<�����0��}�߄�r�)T�I߹`����T�u�ǌuq��S6��j�bo\�V��2�N9_4aMY��v8�teu���ĎH���ֳ�;k�k<��ĉ;��i�r˸�Vt� e�~�W W����*Z�)�詡�2"U9�c�Y����Kd���̮��`�P3��� �E\�Wl�Sn_ �W�]z��f,7<&ɀF���R>s����Ē�q!i�5X��Ǥ��G�L�����׭���6th�1���w|(s\/ԈM~�����X3�'Μ.�/���0�W����%�L��&(����!F$��甧��.���$�K�n��0�������P��FB8�0mN�kdG����@%�sT�D�8�U��a�(k<7�}�Ȕ*�ȹ�aKH���74�	p2���]���6�io�\	����F߽�\f,������[{$����1��&�<	�7$��c�{�&���d��}%b��s��`�꿜�.J�7#��Y����#CL�QEg�5H����C����VS+�v��x$��p�y/�Ȣ1,�z�`Dm�/���H���:��w��vsxʷ6رqp B�	��2�괺KZ�Y�|]pP]0����?f�Kl�;R�_��P�7AI
2E�25,zg�EF��ѿ�Z��� ����r�i�������
�B�� ����u`��dO�h�:Zw�7��^�M_(��e���T��n�E��>��;��,�aU,J'��ɕ�k�#��E���"1���t��z���<ϔ^ڈ��>;����w��ʺ�7�yPxF�dq�:9r���2V���J�M�����li�m��8�A¡�հ5��;C�L-m�^�<H(z�o�瘕H��pjm~E#����Q�Z�$-��Vof#����!�O�"�|��7��228L$c6�mH�E��S ��F,�+.�Yٗ达�Xe�Z!<���L����`�J��I#I�~9��C�qW�H�,��N�`:�f�'}���n��[f�s�C:�ޙݟ� �M,�����we"��(L�¤�5��E��H"3�<LBzJ����?Ұ����.x�䱥�})4C|/�=d�e��*��on�]G�P���2~�l��g�Wu�jNf�45 �Z�I\]p��*~E�<�6�ǔ�:��`x��(�	ԁ.m49�
�ǀȸ53V���b���?L�ϝ�R^�G������14�8w�zg�5��b{�\�� f�f��SI�D��&9U��o������r���*!��%-�7�ÖH�l1�496r��{-�E����"�;I���]_�0|Aɶ��d�H�?FU�%��U�FL���+�W������V"ˬ�{}4V�:�74'���f�<�(FU�¶#�H�ɷ��[EG:^�� �ݼ!2��o'�ƙ?SQ>�pi~�t�qL2s@�Vi�O�w�?�;a0xͶx���d���1�X�*���jl�