��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�#!��{(�N[V��/2:DY��6���T�'��:;�5(8���$��Eʀ%���4e�p�;��a����^JN��Z0����> ����Z�� ���1���C���Ղ���Z⥃^��մ��%���ݎ���
E~�(6���B���$�i�D��%����?f�G���Cy�����J���ǩ��5���z��d�޹��L�t���M���TD��Z��oW�����l�$�+{J�M〮�
�qH�37�t��KN�s�$D�^��E�޵�Bl |$�[�Hʽ�y^I'V7Qt'��ѣ|DA���Im9�-���Ww�qG��>�soҐ*��^h����[��<�Npz�沙�����@�-���\(�fR�i��rDz)�J�}���Tw�ǳ�u��%��	�w(�U\���Z����u���%���9&�c��h��h em��N�(� |���i�L��t�4��b_���A��7�VR��Vr��R=�f��8�%=� ���)6Gu@[��i��U#�ޔ�-OS��Ӊ�v8�'�w�l.7�ʋP<�k�<"W���	2��X˵��
2��0¨��q��	Ы{�P��m�	���%��K�O����[3�;c��D�Q�I�PQ5��,��ձ�{Pb�#����3���51�Պ��EAyl�������xZ��⑞־.x0����[�g�٨=b|���j�|O�<�]��tԠ%��h�����>l$�'RG�a'g�ա�����������N�T�s����a�
�Ȱ�e��Ӳ�����D�9Խ]��}��~�5�p� �U�s/�i�$AW@-5nMĨ�U�P|���Rs�
��k�`%�"o�(�汢�ߎ?ի���tDg�*��3�f��h<9 �,���d�v�0I�KWI���B�(W���[jC�^��b8V;�ů\fAG*���{���fu�Y�$�s�z����$�i\���@�C0��z�@b�	�`�4a��c���%I��a�r�_�v��?���S�H@P�H��ݕ	�y�8�]�O�T*x�x��u�hq�D�l�X���g. �f��!�#��2�V�W���b�L�>��A�V2d�OI�U|��=�$��Mx�/ӳ�^����S�ꘆl@&<��.Tޣp,U�;�xħ�إ"qJT�j��q��,޾��F5�|c��PG�;������b��#T���z�p�%��IR��8_����6Q�`�l���}7*!4�tgU��SM}UB��B�v>�V8�����X���Y�A�o�V��T)e�O!�nB��U�?�qB��ec��HNd�&/T�`���3XHL56�3r+��*�hv/P�N�m��xoPI<���szC�1��?��:�)��G�a�N�gȮ��;�P���a��N���=�Ҽ.�Gi>n�}uH�K9E|�7���[\Ʉ=Yߛ��풼�uZܩo&�&��2���<���=S���Ha�t0����֖�d<;饉��$z�x�Q����>�����ax=�2ۛ�������ޛ��nd�׽��e?��{"ɍ���n�6�[���J���i�$�{�p����WD̃�t�d�"�2>��g�YH���}��(��pa��B����i�E}l��G��x,;�ESm(o��-�f����LEwy�	�*���%ȡ�[���j��TAGn���dno�U�iW�e�#�v�Sۆ~QJ��ƺ �n�]��X��:)H�ǁ�./��WG��:�+GR�q|_Pe���W!�%�/K9f\�A���kr��˚a�s�ge�2�����z�|�Qz������]S:$��K�a����7��4=�-$r�x�12qjg�7���D$M�`��p�p�=���z��a���e^ Q���I�����7	2�]�a�D �g�>���\���_�T)Z}���Z)��&�$���G�L2�G�Fn�/���2q��`�31sRj�,Dw
;��PKv��!��a��)��Q.C�A~�۠3?Y���,]!�d7��|�������`񆁾�T@<�O� b��l~OĮBM�ak�]�E_���x|�:s��}-�-D�ҝ�6"���;�C#ͧ*�!#1-pa��_�;|��s<�,rHq����WЈ�L}"���S����:���J�/2�)����.����w���"��M�k+˭�C��imoS�G[�=Ŝ�EDV��ΐ7��KvcdP�7�ۨ!�
�7��{���}3�_^V:z�N���&��i��#��7&R�k*�X�|�l���>d6� �,0�'Ć�Z&�+:�_�CO��ܞ^5B^]UO`O�G�PH��a�R�t'�|FC	1��yM皵��ڜ6c��I���O�1ٗ�t$�w@�	�V�(_�~���Mʭ)kq
�ͬ��V9���#/�i�h7�[+�ț�d�Ye9��E���1��������9��Vh.�V5�&�{�a`��①LZѺ�8X�s�.&3���
�tP˥py6�W��f�lP&:�d��O�3���TJ�_������G����L,������}@�\���D�o4	vܢ��
�Ż���VN���:�Z�����$���g!��+�҈�Ipl_��x���la�v?D��F�"������tu�C VP>�͌NI����܅>��r�����,s?�4=mT�����h�z��`z4C��.�άZю�/�h���G��/��	����O����K,���-gyQb��;3������M�K@p�L��� ͢h*�E�u#	|��6��BZ�%c���!��ȶ����`��F͈�W�M��*�l�o�'�R�'2�M��4��4=�9D�u����Mf/�G'�'v/3�G����i����!?C�:�wI�?����;f���t�^W2A�����o;���P+4b�{�ı}�x��T�x';��AC͢�C�����V��g�Ό��Д�X��l.u���io��5]}r�#�R��+�K����\�������8�5
LǮ��[�Ъcoj��4G�x8P���`��y�t�`�)����+�=�.���=�8�r�J7*��g��/�uk��O�?���2�T��N���%u&'�T������J,�p:\�{��B�w,Y�Jp0�|�u��7~PL��Mx~�i��q�밓2Q��L��h��N��+��}�8�HhG`�o�i��&aҮ��³FD��2�Z�iδ�>f��;��y^�Ox
�qI���"�0$UK��
�f�B)��D���؇*D��JM�4>R�Bː����މW 2~�B���=��-E
��P-��FM�����g*��&S2�S�6�Bu+��S�)�!��p�ŮSv�h���׻�pQ/<ϧ�p$��Q����:��Y-cO���M��7�:y%�U���J�C��s���>Jc�e3���.�(�^���<3��*�]証�o��Xk"C�T��v���`��q$�"�r�{չ���t���hLA�~���OO';{G�������߀n��:���k��A��e%�|j񝰄�� � t��TɺX��"��Z/6�H��*)0k^}v+��ۃe's�`��(���H��S>��ܧ,��Ըuy��c����Kh��N�oیݕ���-�/6���b5X�a=��p���ֆ�S5�]U��kj�q��z�^)��3[����œWi�oG�S�4�j0�a�{1J��vݥK�\���i��o�s��p?o�Ԇ���d޴�t����,:B�IC��r�4s�+Ҿ|�E2�ա�V��M��+9|�������1�6�Xo\ؿ���I{�¾�K��6e��0��KS�5� 1����FC+��c4�?�k�X��N�f#ғsˣ.�gyirO˞as���`����[ժ���p����<Ҕ*���Y�9@yְ���*��TC'�fi�����������K@O������Ĩ����$R������-�>tiK�~�a��#�}I�����s�n��>q?{��^ŉj'׊�8�55�	'Ab�2����󓂨��{�4ɭ��l�VL�ȇ��2��5�>3����v�3=}�B(��	�u4掟��L�\�є����Y<K�9�kHF�%0F#��=���f�����#C���6�bP7V������Iq�V*l!�-����0Cµ��֝Xc3�j�5�t�M�J��A;reuh��C��?o83��v[�eu(�A�7-o��Zm;I4d3 t�x��I"vc4��(�����M9�?�oJr�T�����b�����������Ju��"8�'͒$ǉ?���UfsTl�2�����4g��u�M��"���R� �+d�}2G���)wk�uJ��k���\��Tjo	�ZEh؃�_f��BQ�L5/^�U��XԪ$ռ_'�I^íT�v�����'Z��6�����p�J��_;��>���	���<�k�$5�B�N5='92�]��,҂��2L
�����8W5�?c@��<ղkj���|z��cu��r�e�@�.�+�X�r��X1�����"L���+� n�(E,[?I�sI.��z�PX���"B��M�ǉ�2#�\�U���}������cs��.�:Y�D��s������[��+S�Y���	��Y�����t�pJ-��C��C��XF<���?f�� �]@Q&y����R��p�3R؈!��$O�xd��[�f�V'l���ׁn�S�{0�I�ҔI�<W/K�Kg����ۨW!%.��L�˵�C%Ѝ͊��:�+�;�s.>�O�������|�Vlʺ����5��$�vB��ohJ�"�J�;ë��J#����K���%+o�?�}Þڣ��.b�~I���պ>5c�]�[�RkP?� �{��z�?��z2{���7\m��v|��Asڗ<��t�Y[�����~�M�\-a���̻�H2Y[C����Ҿ6���u�����iWX���Ӭ�r3�AG ����0����L[A%	y��� C�l�K	�ڊ�ͷG�h}9� �&t����F8(gN�:AB-o9�@���Na \:x���T�Vr�l_ՑB7�o>B=p.0�~�NO��@WP�`����&���/
��=�p��!��,BI�k�	�^wWF����C��2�-e9(��N��m˪erd"���jC����{ I��j�^�Y��r7�T�<�I'��P!"Q�E5��՞�i�,5�z�!�����T���S��+\���	'mg �=�5}}�V
�}y�����2�|q��<0�	%�_Cx#	s�F���6��<?y�&gׯY���r=�5c��"�0������-��Ol
B�(�}��'�~_y�1�&�-4�&m�%r��T�(b`wMUy�ng8���2�Lݫ_Uj�=�pGI�+j{Ǫ��eO`/!�0�(=��*BQT9�x*'53�ߌ�y�l��:T�t[�[7q����?�|t�7��˛m- ���@I]WqH��ٚ��w�S�-��Ƙ��ϑ%�&$AQ'%~@`�~��$����f,�o;������R�x�J��E�s}��S���R"м�ʣ1�n;��3B�������Y��0e�2���l(`[,�-U�D�(!{��&���pF�!)H*�#���Q{��GB�-��[�\�h�C|��UW}[[�x0x��8r����%�����j0!�[����K5�7���x!��û��60Zq��G�����K�3u�:7`�]Bf>������Y����)"7���ѷA�C���1M's�~^����<]hpU��F��(,�B�c0O�C�eY������C�����=�LW�og���Br
��3/d�P[@f[{0�b��6�d��1�	3�.r3{X��-ƽ4����6�ey]��k&}*5��cKz��{z
h��n@�)�8d/�YTb ��x����T�q�	 EV���^Z�*Ä�s�t�&N�ɯ��jG��z���6ŕ��z�j �1�P�hi����fY�.�S���#|��N��7�߲�~m`�����
|�Qd�7�-�vO���k���Z�,�C-?�Ft
ɿ]���uW9�;��/T����WY�kRObi���ʚU�����Lg/<l �m�1�σ���W>~��gQ�:<n�%�ԁOt�Q��8p�h�L��3X�5R]VI�ŨB�5�@;���qhkɪ���Od���B�����M?g���Kq���X�,[���W�����7z&�Oc]�*"rL��+ŧ�p���^u���y̯�I}�ל�۪�9���p���<52#�Y�h�W!�X>�t��D��VR���e�[��^�#���H���S�@Uf��v!|�$��%������=���&�u�(�:Y�}�W=Xw�ݛUpq�ʻ�Jp���ߏ�(���ut;͓�\:�T��q�;�� T�Bt�Q �sY;Da���8�ĩ�TY�)]���������g���\i�;b�JEm��6_��a:ᑆS�{���j�j԰>��˜'�D���V�&5�x�H|#ch���6f���_
�V���.u۶���#�WA�R)��Pa�-��{���S0�����_�\3�@v���NC;�h�V^��B����7��8#_>��w���/�1�:��։x���g�B��ZI��Q��J�q���;��t��}*�tR��$������I)���J��kh'8p��o]Te���Pa���S�ar<!̺��}{�YHq�� ��X��7��#o(
k̿T��Qvk�t�zTy����pYŐq*�'����z=�؏cLu��A\ݖ�E!�:k�O���<P���c�c9��͘R���H30y���و[oF�=�N ��"1N,4�2�"���ύC;���@����ҁ�r۩d�;��*]�R�8i[�#cp�,�� @��jω��R��	�iq�."JM���ˮ����=skq{_F�Yg����5��y����"��uiq�Ϗ�X���v���+``UX����g��*�Bj��c�wՑ14+�W8�f�0o���� N��r��.�w��r�v�;���9j��S3�P��F���{��>T�,�!���>��Z�k]�5��*��^#n~��l�|A�X�o�>\Ć9h�!*�[�s�@���fN��@k_w���gRՓڿ��Xo�Ѱ������|�f�<k������
�&�T�.��݆4�ڊ6o��uX��:����