��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^�}����}����'�����U��܃�Je؝b&##O)ʴf2���:e!7��;�C,^:����C3����{�Eؓ�E}���	7�`6 �e�&���7ۺ���͒PA%��� q�K���\��Ɂ����;D»QY|隷�F���e�0��j��)���[A�%�� ��I0��T�?�ޤ'k��[�W�����?�{���&Tɍ����7��4�Ɛ4�����Hdo+��Ch�nE.��MTόV�	��1̈́z=�����^iKӈFD7�"<�3.ab8���r8n�X��}bB���+����B!̦�`���rЩ^��㡛D��Z9�@�v^�$���G��Ѱٸi³�Z<�j���v3������Z���%LTw���z,�2\/ʏ����y�>��T��k�a]W�C�Sg���� ΢�?{�hI�Oьn������{�&�εn�
U�c����s&:�No4B}��P�Q��+�H�%��?���Ev	I#��jvO���WOPP^�nh(�����7�坖|Y��{g4��&�n���I�?��;�h��t#Z����:��q���g�z�Ԓ���@����n T96��ΰ����ɹ��@� ���3�S�yC흸�� F��|��j�{��nN�$-�@G�#��a�]��֐���aU(�k�?�=�u��
L�!$��Skن1�
��ޯ�D��~��CP�� n�����~c��@��u��G��tբ�S��{�Bˬ�j�v���څG�W��=,PNGK-�^�Z`��`T؇�k����YGO)�A$\�5�2�K�9zr; �����s��`�%4��2ģ�c�\����l�w��'}���?�2g��cPoT�	�����plr����F���P���������ˌ ۛ��]
A:�8�+�D5G>dU�߹��}���Y�?0��vcF0 F�h��?�����!s����#�U�^5���8|�������D��g/m>?D� %���������%v������5�u��V���nN�9����1y���j���b	�w�y~�	�?�SƂys�}��B���A��vM�4�k��������p!ߨo��{�eX7�|���x񛁤S�6���]�M����]λ׳-�=���vș����^ /D I[�:�!s�	#_�zW"������Eb�7���"$��!���:��A��)�8��u)�.[<��9[�p#"�>�G .U�T�E��7؊~$��5A`��6dj�Q-0xrUr���WT酁���I��:c�u��(�ϗɁ�Yq[VF�ϗy��#��3��dz�^?v�s��#p�<XI牡ݽ�K�W4���ˊ��J���J
Ps�7(:�5W�ܵc��i �0@g�a�������Wސ|��y}���X�7�ޛR#�����9}�p���΁���Ӥ�
�^`ž]"O2E�_##g������/�=��:��;x����|���L\��W̼8M�du�����*���.*���X�s�&���؏-�:���3����I��nRy-�T9�Ju����r~F�j9ܖ�U"E+�}U�νU��t	X�zͺ�A8y8�'�4�f��C��b8�[����.�mq�T�wZ��;̩��ȧ���}�2`$����?>r��SL�.~z���K���1r�`�]���w{_�KT���l㣜�""Z�]\���ϔ>M������E�1��k�I�	���ɑ�Ϳ�ǙjZ0�vٚ>MC",|MX�D��T���ɶԦE����MK�E�{��2�b�����p$�F��;d�e9�}�z��hVj[m7�@�4|�����M��B8���iKˌ�
���|��p]�-g���0z>N��)���,�B�I��s/�2�CL�i�|��E��3CW�_�S��I=R��H�3]d��VXn�T@p�3��� �Mnt����S���������%��- ��� ��82����8	ͩ>�1:�c=@�H:�+�R�%
�j���oE)R�?`�<W0��)�A
�a1F�n�xK���F亂�bT�&;�a�ށU����
�K�V囮�-� ��t�d��su��P�.ϴ�"�����ᓯ��p~�J���o�i��a<�q������X��ٹ^����C�F�k�Qh5�\{�����%'�H�|%��W}Ow�lHI.Hd�HCeX�#�}9R"�)S94�G�M˰�î�ュ�?��6�lґ-�E8�%ܹ�3��#T9��F�	ɲ���TX�?TP?؀���o0d�Y��xd�&[���}p��~rAg ~�RU�uF:��ܙ��	�aa�+������Cg�jXU��ԓ9�xG%D�`��h��k.�-��y�k&�=����0k���є�&g��Q��Ca��ͽ�O���"� �����B�^'��y�i�r�SN���v�X`���$zFXx���! �'�(��6ҳ�l9\��+�;��3U�<��X"��M���+Q09;�����5L*k%����p� �����z�����P]�x_Ī~,Q��������딙�A��~ySpDa��iٹ�$�\��o �	���6�O��O�W:�J�Ti�g?�jIGΛԦ�w���4"	��Pk�������Rr����=k!X"mC�i"�H�V:̠��%�T�RĶTF��^؏( ���~g��؀�vk&�W�\<Q��dnyB7ϊ5Ms�ъ�WXX���~.��N�D�.F�h� ��K���X�P�"ΐ������2����l��4MP�5o��fՒ��	��=]�������,����LN/#P58(&I��SV����K�t	o�a�"��V�M�2�r�}���\!J*���}ae�Z���cy	����1ʽu�ݘ
��r���#x�T�O���V�\iB���;�������h�S<��͠ȁ�a�n#u�7'��f�D� T�1��*��^!p_��:���Q"%��'�=.w�kfiB�<���|A�;8� �����߼�#�'%U��pQ�T7�Cf|�R�Dƈ�*�p۱�xC{�&e��i���w(-
���iF�B{� _�7Los2ƍ�Bg�m�'I�}�V3���L�AX��1��/Ĺ�c����7���dOsP�m �~���W~��T2��ْ>�V?��jU��e��K�����	� ��Q�M�Wuq��e����D��Q�ءE' +�V`�b��7W>I.���Q�S��:d����+]���Ù}Z��A�q��	��S롔��% Moڜũˉ�¬:�ֱb1�IJM]e��w^������Uä�γw�e�	������2��T���	�	
*)H)Onp���LEk��,���\�w�&�+�_ O�з��0��i�m���އ���0TI~�I������o(k�>(�P��ٔk��H_�*aS����Dol������-E��q��<�n�S���_#���8~��sw��>������j�R.���J�[������&�1��.�^��	�������Ch��WJ��<z
VP�{�V�"��+�6zom���(�uZ�.<{�s`��9��e6Ȱm�ٛ�p����ىX����w{W�l�6@3(ڣz���Q��s�l�&<�.w,4[�4�T+}hZks��2�$���ؠ5�Z:��e�(������X��B����dD�nO����4������GĜ�e��<�,`Rm�ӗ�Ut�����B&o%B���l�(��W\�rJ�}E����UY��S���)/x�t�T�*d㭏]�̵���HK�#X�D�	!ǹ�`j�v��6��O�IV �D��	1�!�.%�j��X|�H-�p[i��d��!�y���u����nk� �5�B3���+Y����QE�������!���s��a�7�|�S��à�)�=����P�_9K��X�{DV��h ZOQ��'�2�y�������os����řz];2@Ɯñ��S�߉�Ӊ��FG����m��.4tY�n�wk� ���l�~8yVM1��P8�������4�]G�]\xU�O��	߰����Ҧ��bP�������qÞ�{�-��5]��
RFח�?��KutrG	 -��f�a\�To��N�����\���-G�k�>����U*j����+*Ӛ�+�ζ��/�*�F`��0$"`��=�W>�xTN�ˋ��"3WU�w=�(�v�$���p0(��W;��QI`����k�)⋗��3J��.Sf���Vb`�k���T���S�
����IռXR��6im��_�j`�
1�?����Aa�Q�A3�܃$�E����=۩�{��+T�>35����J��-����{��M��qW8�&�^Qb��w����h��S�e����V���p˒�}A��(4����R/@�0$�|�s��(aHv�����,eY9�=�~�h�ɚ�����t��\�����J�09����9���W���q� o��؉3d^�i*P�{�J���G�� �S��u� ��f-ߤ.��eqP��ed������	5ф?B���6��6�6�F���ir�'Pt~�A�T�q����J���2��ډ��n��*�ntq�Y40X��̞����Xt�?.]i����J?�w]�A�l��xe�:�������fG��\;[J�I�nI�u�W���u�z�> �۾���D)�)k�"s0����-��(�Fၷ(��彊ێ�Y'�M�u�W�u#~D�V��y���ic ��)�N��J]���rE~��o���1�j|��Q|�"R��j��4���;����?Q��O�<֍�4$�I�����T����P_�y���ҳ �������>ӡq�E�.]Y�������b�T�[s�zx�Sj��]'�Lu�,��� ��VB�^韧ѩ!�*���SVq�ۼ���-v����`�}'�3e���H�MTI�/���D�����?q*&\$�@�C�2�~����
�%���i�CP�8�&2�W�O.Q}�g��@{�n���?&����佗��vJn/	�0�,���Di����6��J��7�J��gs��,��DS�)�v:�"�4�]m�Ud�#�z�2�#u�X$����ڜe�g��rd���54Q�|���h�Db��7���j�u��We��'.�Y�R�w[��-ah��}��0���p�����ѵ�D_F�����iT��c��C�O��*,4��5G�w�)��Ī0u���1�	�KW]��r�Cl�ueB��J�d�p�,��]��r :��H���D�߉i�y���q��HV>!k|�~��3���k�Բv\�����Ɓ������",}�%��P��F!�֢ɾn��ϣ�;���xM\�t'���XM��u;g�U�&�P ���oj7n������g��Ѕ�Lt����8� 4����CcqQ����H����q������}ֱ���u���k�K{��?�{
�A���ʨ�����-ֽ�72>�t�H�.�c��TSl(.	ٴ�����~��쩙��F�%zފDiV��[�g�5�p��#�ވ�A��t�NF=�Z�fV��f�B@�jc����7L,tWO���H�)�Y�;@�r�x R=�H��n�#�1�Ж�?@���H���Y̠@%>��S�taƩ�����Nd��[� �'��uf�� �i�ߊzP�T'*�lR};���fS�c}�5d���>���D��Dӣ��F蘃a���'�֨l�h'���O��
��uJ��ۻ��;h~�Qowp��C��5�`W��$	ykj�w]�19ȡ>*�+�9���T��p�l Wv�Z20r\���`^��@�vl�mn<C'�)���q���;�GBd;H/|T;q�Z�Z��5�/�E0D{âڹ��W
�w�v����IF۝�-�%���~S=}F@���J��ڽ/�/�#'jӵ���A����^ݧ�`:���a�f���}��C�hM���"���HYx��T^�OS�)ɘ�_>���2eP�����솘�+�q$~/x0] �[�ZH)Ƒ]����e����Y��Rt�l%�
�>`S�ڍ�(f�jZ����7ܲ�0�{�:KVyhl��LՐ@|�0e�"��⌟l�L��U�6uC��F2��q��!�Á-��N�!Ŷ����`Ob�)Js[H{w�a�GW���E�s��mB�N����9^�Q�Ăp����������Q|�J+IjJETn)$�Iz��d1�ߢ��Y�����VExg;��-7ɰ�����Y�����s��^!����y422ы�=��D�Ԏ�8��@q�}�R֕��Hfз�0�q%
�o���F�?�:�����\��Pc�%+7x0������R��-ٱ�%�P�ѣ!�3x5���ة3�O�#|c�����~g��)d���y�Os;Z$����YQQw�c�>/����%�K<Up.��lǾC����߇�����Ɠ�pY��8B�l���� <�ݯ���L����A�<*VWo;��$^&R�s(�de"�t&<?o�h����;���L}�7}8�i��cu���HVWf�����9�I]�ӮR�\b_�w�:M��N�dT��<�t%� O��S|���]p���W%��m�ڑ��l6A@P���<8�,ȇ�A6�>�摢t�*<_���bP6�iXcZ(@���U�����q�'���0�{b*�1>�jy��$X
IHu�v�@4��P�Lb��oo�)s��UM(�W�&��^G��4�G̇B�u, +�tG>\��s�=&kh���>��9w"��|O�r;�Һ��QQ��r�2[*�w;`���5���Mr�QP��-JIT�: Tk��ԞZu= M���W�s<�5C�Q��A���Wx2��bw���'��Tq{�]Vg/\5��Һ#&s�����tro16�]���C��f�]%�#�_�4U�B9�ei�	����a+��q���o�W�D၂5g��=����1�ѯTS�?��mv��C~i����):����!Wh7YeT7�m�B;��0�C1�f�шg��OVT�#	��T����fJ��m��&�1-��Ww�m��ΰ81�]�e��H�(�1P
+|P)t�O�I�ޤ����V댱�.�{dA	�YP��}�������'����$o�Т[���)S�i6�H^��*���6�rz&������mr�xJ6n��И������UY�H2��Fm.��وm�֜�3R+����,醦,�;5�8a�
��BUνdY��vR�K=�iX�Mf��*E�zI<p�ꕴ���kl�F	@�����Y�"��X
�f�A��Y��l������br ِ�Uf�)���\�ܨS|��)"MA~��tc3h�X�UEM��BT��8��D��:[\�ng����U_$�� �$ㄅ���mm����b�ҵ#D�Ueh�/i�E�{�yV5H*;�bXS��Y�I<�O��z:E����'��ZϹ������;>
L8��'(�	dlD�d��D �%C��f���r�ypk�����*�@��R�����a̺��G ���3T���y����p%|Cͩ*`��:�X�I�@���{Y������]7Ѹ����kڐ:�	����R���i}�1���=l�,Ȟ��އ"�j��f���s�a�NSPq2�.9R�"�5tvv�_�vq��x��~����3��-8f�krJ[�b����Jas�7��KX��$밞m�S77��}���A�L�,��� s�ӷ�l����ȿ���
��Mwڡ3E�*��p�T��pn��.�ɧk��/���|ދ�CH����B;R�����u�T���5�����@|������L���(�V<;~r�;$Z�"ao$�>(����q
�a6�9?R:l/+1���_�p�GI
(�0�n�Ƣ��W���k$�#F�h��_F���֎'���4�`hs�.�(ڳK�|�#;��yy�����tѯ�d�T� 0���k�xI�S�qm���8�+��ջ��b�'�B��D:��:G�u��r����6��q hY��^q�,*//M�1Kd��<�J�}jL#"�sA9��p&�-�d��!�*��&�3��]���)�j�vu�y[) >N���3] ���6݄��*�Y��	j��0�p��O�M��|�Q��4_ݩUH
�]��Թ�5 ��nZ4������}�ͫtr�_�����ҕ�]�țmHc�/�.��RO�#?��2n�X�C�v�6��>_ѤB�1����lٝ��PNJ�9-�p"bo9`�Bz�n#V��f�@�5�k��~,��?j��R�V��8!�܀qA)��-�v�ɀf�l�Qu�N� ���2��B/Q�k���q�1�zwȟ{��]#y���e^�`�-�]݈
�v���'ff��݋��:�9���u@��ţ�a( ��C���uρ��>*��|}�6Tf2���qx������\�8?R5�.����t`�(� <Ꮔ0�B���HA���S:�НD��\[��=������[XNs�T���:��<FĿy�\��W�MSJ�5�.�����#�Q7���ƧW�I6`��_�W����5�Q�n7�Ǯvb���_��0m�Y�P�	�Uw
�K�5	��N� f�普:�?�9�ǆ�1�įd�Ze$2��U���>z�]��HPn\���r�T�Y��<�L�U���m�{��OX���1K�Q�t�oo=;���lԷ�q���<�h�;���ŭ�G����������Q�Z+x��.��O�h���>Xe?~��e�a������lh�������MC`�/5>fQ@��O�������Ȁ8�J�KRW�� 뫜լ�FU5��5����k7
�����i�p'���Av�!aT���V����33+�R�H�]���,H��0J���wv����ln��ٖ��X��TB��>�m�D�Y����n�|���
� ٽ�{)w�/�\9�,�K��np'55��S�!~�n|R�y��h۲� k�R�W� �%�l�6����0�H��uj�٢K��OY��c��� ��H��s��7|�_�bON�9&�ٽ�T�0:+#��fj��.�
�ۮ�kנP�e�ȏ�BgB�\���y���e��{�1WZ"�2g�/%����QE����gR��?�(���	&��� 6�)f�R��w��N�J��Ĵ" 6H�UJ�m2�5�WY����*�k�hI��$+�O|C�yB.%^˴M�� [�i���+�}JT���x�ڠuǶ�A����x��I�>��.�r�#[�>�|��#~��Qc���]cK��f\].8IkE��b8�A����1�ĳ��1��^醓RAX�A}��^�D��N����ǂVuHS��p�ma����w#��Y�c�v�A5֥�c�"�ېbuOB��~r��1��g�������1E�	 ���>���XW���|HWDA+C�������]��I���;��;��� ��3@�:�Z�ٺ$XKE�5�����_�_�q�^�6�m^�F��|k��n�HQ��^e�]��~N4��V�}Ac��c'*������I�z/���;����(䋻~���9A4���R�Q �+h��o�z�m�����-�Ȱ$=�w�ֿy�p��4���-�ˢ�����٭<Ξ��ތ�e�wa�
�c�����������=N��ѳ�|���)���
�:#�����'s��V(%"jt��Kk�cn�~�M��Y�\����k�XT��al�+�#?��#�@����)�!��T��IjqD�]Y��u��Q\����>�T�D�I���m�u�[����J�VR�uO/�F�rڡ8&�����T��k5�&M�o4�Cg�
WoSPܞE1���f�G���h�� �����M�/�W�������v���>�Y��~@��������m�	^y�����h@4����X���V}G���l꓎��{bG��Р"�h��04�%��u@�- z�ϟo�܉� x0]�_~����0�����n�-�n��e7�/���?Uׂ����79�?��=���K����wl�#~bR����	��x͌�D��e�v/X8�Y����Q)oM�c����^@�~�Y�m)��->�+d";+%����.�N#Ak�W�$:��P���'���!ؿ��=
Zv�+v�t$@^&�����,�̓<2�{��tֵs�cO7KS'��"�H2��O�3� �\�l��#޺�F�}Ԇ��2���[��~f��ųbr#2��ùD�x-��P$s�?^?d^Q�:=4A	�}h:���?��٧��x��o	�KD3o`meW�2�sA"E���B��q\en�D_�oIœlǓ '�ء`q��w$lf	�c���XK�n�:��[�>p5�;�fkd���Q|�:̛����n ��R��̔ֵ�R�T�|�㼪0����ʿUA��"2��SCG�_���3G����П-N�}�õѭ�����󋟗�cB�N��||L���ݺn�x�j�3Kb�J^����^m��/�� Wz1=�m�SM$�68P��u��q<*!�J�9���/z����!bL��=v\<��1q���u7��JL�[�W��Z��Jʸ[����⊚q����g;ob7�*c�6�Cp���G�8��TI{enU����ܳ��vn�ɋ�B�������I<rm<�0Fom��lZ�L�%t䜋��ݰ��?�B�5/�y8�ӽ��V���nm^>�O�j}"�s��u�
���L� M<�j����R��ܞ6���'ZK��f�E��f�,HE/{Ԛ״1(Tغ_ i�o�����0��-(�������-��(
N�Y�>�j��5��2N��X���E��W�]E `lp��."�1��{[���>}��e}���j.�FB�*+�SW~�<'M�����T�y,GS���Bq��g��{o�h�E�RzP���M�vM�,w8��˿=G�ks�e��Lb���Qo|�F&�A_��Vk�WV�wxK���)� ����z�����Rmp"�g�4`�C��Z���"�u���J�pH�b|���Oj��������ܤ]��a$/A��ߔ���N��Z��Q�Uxη^�����sa$if��_�?�Y'�6��S--�,�A���Ya�=�m��j�1��{:l�R��(�� &����4�M�p}�r��C�x�����i���T��:��t�3���8�-�kH���J�n�<_-�P7t�.���֙�����=4��J��FV�b(���H�7d� +��XL�M2*�t:��`'�3։Ȭ�d6I
�T����IDS˔����XU�軾��y�n[5K���N�{�J����3�l�v&�X��)�0:"�ѵ�1_��F�M�9q��道LU�����0v����2U�&q��U�s�Ԭ�3�v�+���t�ϵT��%����I�ߙ�7��PP2���r	6D�7��X�x��w0w��_A7զb��l^�;q�����e�%������Nc {����J�N��(<g��I�y�n2ۇL�Mo9\i�3�DH�S��U��$SM%Z�zEG���q�I)�t�E��2��y��e�݅IR$lk5f�aN��pnO�I�L��])_�S�@\�рӡ��'���0��±OQ�������O�`�O��|����6�I{���k������0�f>�T���	�2�;^�-kU���[n�D3�B�o�A�ZT�?�TO��q7\+��.w��{	ѳ*H-���$�\%N%h2�ّ1�gː��k��5�r���� ���2�6�8��"i��(�g4�nK��ֳ������ghN��,(�@O��2%.8�K[^ �)���V�{ͣK"_{����R�k/�}����z�R5�\0�:J��(e:5;c?Ů%��k�ȝzZ��\,�}qm�b��S%�[_�TN�l�Ml�<��%y��aE��yٜ����q�\��D3F�����Cb�Mb_�.��AU�Ò��rg�!4�����*2K+}�K!{?KE�����t�\pHA�f�(��]Fde�ѴА�v���o�v���:�o��f�Ԁ+i2RPg5�|Ro��B �r�u� \��Q]6��#Rӈ��*���,$�p�c�*�7`�Rw��|"'�>�4�(�l�j����c��4�|��8�]�|�2��]G���8k�gH��!uy�5=z}:JH��p���\ �e�O�����q��w@s�A(�Ws���>6����7�\����R����|���(�̟�,qYR�
�l���"�"ˎ�é9�o��_Ջ䙲�.T�#�4�c�Kϗ!�0Ox�b͠W7�Ӯ��Nlk^į�YL%���'@a�B3��r��Su�	�#���T'ɟ�sm8���5*�Y�(��7-��t�u�["����q/ĕ�j%�v��)����`�7�tHc��Pr'mWp��D��+a�s6ؔ	a�I3�(	RW�@�����hdU�D�L��~��{Ք@�k�6ʮ9���2/���	ܙ䯱�Y�{u����dy�K�����U��P��E��4��6�M}�=� 5�%�Eː�q��!��t,lR~�3�m�fwmJ�M�X���w�%,�	ʕ�Jg,,s'����<"���E�:��6��U��'EUðf:7�w�j�Ǭo�AHXS>9�Թh�5�M�/�&�Zr�4����J��cI|l���F����0/�Hճ��!�s�0i9$���C)q��2���\ӡ+ί�9G��RzAţ�k )�A�_c������	��!f��3�<٠�͡��2'� �x��>��G��n���!E�ȥ:n�}	T�����N	���-��evK��� C���	���s��A�A��-��萓H6@���u���AvD� xP���+��$x2�yq�ҳ<�/�L������klH	f��K�l(f��#|�H��ՙ���*ᾴ�O�j�v��N/�L�:7٠B���C�M�������3�%tc�%�P�w@b�OOe�19�d�m��
&�	�_^Mx��H��ˬ��kJ��a	�V艨�����T@�#���,���@��cT]�ʓ7o��-�ޯ����^h¿��v�"i��z�
���t��	�� ���>4饖��[������ʪ5PFj�Ϝ���m��D!��~�^[��G[oҬ�V��	�1xk3���%a�^�ut�l�:`
T�yKxݏ�{�s:�[M���Ry{�Y��YY?��&>��:G�=
c�Wb�N���a�}��ޢ���x[�Cn!�1A]h9[fa>"���J� yb-��г�I�/�k}�Jg�wS��e��p]0��N�����c���7��
t���qT7Χ�O��_q���Ծ���Uϫ+3*���h}q��3��0ڥVMV(ҥ��k�x[��s�;8@��G���
��x���Gqɥ$�(�$�|�a��w�yiޟ����On��yW���ǕΧ[��&������r�g)$Q�7Mc(��~�IA��:��j�@�ŉN3��Ԃ���0��>������'�Z��mN�y�M�E�Ҍ���җa�@��aLWc�"�$a�k$�ee�[[4t�K���e�o�o&S�F�9��0���qtp��_uy�!�+��bW8����Ű;X1tT�Q���[2G#o��r����{-�QFj\�Z	.��5�F����(
G��Q��2ηK'ڰe���ei͑�Y��'���Q��H|J�}��*]r��*Z��(Ю���������*�.ڋAf�%�o[��2}��L��?p���F�P�9;0�sq�����=x8�;�g���.\��ݢ�bޭW�O���s�>S�z����Dy�+s&K:ܩ �n���;9���7t�30 *�YPG[cNEHQ�vp�s�u;�E#�p'�)3�gG�����&��b�4����[ۍ�<4+a8�!��T�"��.<�/��\B�Ai^�+�N�E^w���+w2|k�B$Q d	N�3�qۧ_;���c��.�帽�H�$%��o��A�Z�Zڗ�g��\��Ն���U�4�c�s��)���Y����+��2���L�0~���v�9t���L�)b�3(V3��چa|�i�5����j"p��dɪ�������q�}l�q���c��r�5�/����Z��؃��:���И07AU菵n�NhSc�U��c Med�M���<+f+�5�S\'��s��Sޜ޻��k^6��BUU�>ZA볶ih6b�8�[���YO��؞�/S�kI�O��kM������"�����[��P{d[0��7�U�����(.liNU�� �kX\j�</i@�����n1���?�r�m�[aO�ѭ,԰�x�&�h'[��_�v+#��X����$I�:ɉ3$IvE>�*��&��*�hC��@q�&}����h�5=>��������&��� ���p������V@����Ur�U�7}���=�FH&Pr �m�)b�1�r�5�����%����^����ӫV�����cC�����c���I��:&��&���[Q�$�S����P��b��(�v�9��CLA�G���t��U' ��{��R0il�����|~��P	���Yģ������S��GQ��$�x]RI�A���?�,k�ݳ0,յ�Ӧ��~��*`j�®�v��B=���%Έ��� BMi��VP�"��汹�:���o z
@������ȿ�:6��|T��f���^�/�r��q��h��S��#�;9S�f�P_�3�������aW���+m��W��Y#Af_�i'AM���tԧ�sB��=��>�):BU}�MsO���R��B�V(�����/�,k{�U�@�8�R�P5S��v��:��!I�Ia'#X�ѫ'}�?~��A���klE�������b�ڠ���ҮӬ{ g�YaS�?`r��;��tU�RR�[48��s��ޝ��J��wjE�(1Y=��>b��:n�pf$�U~�|��VJ�*%�Qٙ�Oh��if�A�!���&�߾�%y�˥���mپ��~s����6���y"���՛�Cb�$�Uݶ�y����B���G$>i	����!R�������
ߑ�O,����T��|J2_��=����%�����&dA���2��1�].*�9F�s�=_,ʴET^{pc�����gOL�P�2��{�ٚ ����,,�j��d��ʚ��t7�[��j@]���8� t�y�hp�[�H{&�B�����W9;� a�n���fZ�k��w_�>��An��ǎܽ���B�S�Ӹ�4Xf�C<����_1��h0~n�v��o��Z�r�t,{��׎S7�?���H�J.��"��G��G�~b;@�۰�tC�u�ɀ�R�R��hC������ʞ�ô��_K;
?i1���㈪�Sf�� �����0���v��9����YL,����L�������a�kq2���âɀ�9�,�ͪ����b��Q�vк3L�pG�6)�{mH�>���!;ȈT0Ӣ�{��(Ӫ�48��@&��3QLUg�����6�m���b�����a�����=r
���"8�������fr�3�\�����֯�e ���V�yL���b�p�]m�n�"�7Ȼm��9��b�-��{�F[^X�ަC~+j)�5F�TР��`�O���1��/ I1�&�DWq�����px%�o�����{��?���3��%����_4�Y�,������Є��-�4ڡ�#���ca�ŐE/k��1<�%�8I(�'�����!*�rfux��T��Gu=���-�a'�7$Ǫa�h��p�*�Y�j@�����q�ʀ�K��VX;��ϭn���ȒA��&��osX�H Bp�J}�R��L���8�sm�*�WX�o�u%��p)���ur����1�nLN'T��G^��s\�T�T@���=u:�����O<�i��p���כp�b�� $J�(=��0� <��^j��S��=�z8���rzq��3�y�0��zC�LW��o�x�fKԁ���t�r�wb[���rF�ɼCb�ݓY�A2�M�#-L\~s7��٦��[}�3�Z)|�(����,���_�!���%���(cӲ{i΄k]CR_D��{����Y30���_�re-o�Mu����eu�(=&��*�i"����~���@�3WD����1�c�S�)Mp�=v[![>�
��̔���B�uY<�N�j�q�l�,��$������0��2���U�!�q���\�$��t��j��.B�(���;;�3w�.��pB��=�`��6MO��]aԫ?�F�.�ho �fʵ��\q�M&����+�!�Ք� �@�rbjY#y��";j��n�m����V�T�B�B�e���	����:�;�L��7џٛ���$�����������|$�}u��3GL�1q8�c/�\*��a@�
�s/^>�Ҁ�4�s"8I媯�^���^)�5��\y�	 k�z�D�mՋ5��h��g"�\�C{�xή�)�aG����D��R"�� �hBƻ^|{8�(�C�$��5��>kn�i��qԬ�����BPJ���[��I�P�Yℊy�烈񕨨#.:�V_����"@/�wX�/�L͞��B��0(���s��g�4�a�O+���C�̒zLH���nh4��Ẏ>M��n����S�"�u�%8D�l(9�����iAJc�2�7��{�ȟCW��s��O]f9;g!�q]J�ρX8x�ë�?,(T)�S��ť��;5��a`��S3O8�7ػ����L����<v�Q�4A�W�^�pi��Β^�h�"�Ǥ�< r	���6���oR�>$(K�)L��+0���?hHK���~ًj˼|��_���S�Ǩ7�M�~��x�a�30]��%���$(���k��)�~ �4�;�?7��*�Pe�5�&���g\�Ԝ >C��Y���rQKv ,������q��EJ��KfjA_$�E��~݁/�����C�҅b��4BY�*C���B��<��`9�31��L"�1?�[�h��bA���Fz�(X?�ebR,;�e�(���$�pz�Aj-���ɗ�.u��3���ڧ��\��"��#���N�=�!П=(�B�S�F��/�V�7�0+'9�(�z�5�KKU[������*gP3Z�,y�7 ��u:JW��b�� ���*x�ˠ�P@����#��1�r_t��w��凙��psi��OIoq�L�(�Y�C�^t�A!w8���(���ɑ^���rʋ���Q"��&�6Z�}�qXM��:`�����╗�S��辸Έ��jUfr__,�f�����l5�&G�Q��z�p��5�d>�Z?��L�!R��&��1��Ń`�*��2U��g����`&G�l�OK�����4	;z�� �P���`8���\߲M�������d�v�B6�pX+"�C��#ď���^�m�J��*����hNja�~\Oq��!��=� �,�wJ���rԇ]p�R�,�]�]��7g=a���ZV�\�9�ś�=�j�B��&.���B���Q�gNw-��X[��.z��xMGk"��a�ͣ�/��r��W�^!��Q�z���4�x��ݘ]3����:O�Q���k{c��dv��BkA��-'>w��k�WN�?b��d�*�o��
r���RL�
u�
#H;�&:x�:+�u\J:�"��g��&���$�Z�,�J�N�w�ڥ/���0�)&�A���>]x'Sx�����U\Ez��/of�*�i` .PƊ@?���8��7��@ZT�<��q;��0\'(��lV��&�=�"�͕e�Z������uڅ�i5{��wl� ?<�W!f��ꂐ�7����0�v9f	tU����ze����";�$K�DDO��P���ְ���j��:�In�����7d�ť�g�'�{��5\�-$�Q���ae�:+q��h)Efh"���ClҿhԿ	9O�ŉo�Ѯ}��:n�H1,
D���No<��2;�2l��F�v���؜S����	�`�+P��i�4E�J/r�.$eR�:c�xN�r��pq=�[���+����A��0Ply��o�b��U�l)�������bqJV�6����PH��S_�p��*��!H����^�����L�p&�}�u�`H��l��_��=��.�L��n(�}��}�����V�K���*��(�\E�GE�F�}ܔ�x�@p(l�I����ّ�Kvd��=!q���2lB18l� �ھ�߿�;�x9o�`.������cK���5KX��%C6���a'}�^��|����$]�X���eI�`p��:U,� ��0��C6PA.$g�qA
�N�Ռv�J���{0�U��L�=�;[�O�1B��^�$��`��b��b�&�tC��=�r��zr��SW׌�צ*��[d�����Ỵ��:z��8q
�X�����Һ�h���%{��o�C�{R�����? �]��ĵ�r�&XQ���"�w�]9��i1���2+1��]�'X����܃oH��4�Se��c��ޔ�L�`�?x���|yC�@�\-��S:�ԥ�_�]�0�F=,�_8㮸��!��ݗ�ؙƃ�HRU%��cp�cyIѥ?�ϻ4wb*�?Џ�ZE�ǩ��u���kD�V�A~�=����r��砶H�&�V��pΈ��\����~E<H�y:<��������맡��#�k����yИ�c2z��2%������3fC�3�%��Xm���?�с�|Q&�,\\�V�^ha���wEG!�T�ԉ�[Z��j���g��#,٠ا?/WN�}�bI8��z�(9���&P���'&��Ȋ-��T
��Y�4%F�B��#�r<�#��(
�V���O��|�!�b4%�L��Nϼ�%�)Z��m@Jc�lZ$y��z2
��]�q'g�y˱u���DJ��ܮ�@�X��y��c3�aOm�j�uڰq��lۛx�~���D�U�4´!�;6��̩�9��H�¤����>q7/U�6G}�����b�w7&K%���(��z*c��lRm���z|/�gE&�1?6x��I	Qtq�2\�鱇�������F���3s?5�Ih�T�������ؠ ��8K�]���e�2m����_�Hj���?
�>����ܻG���먍JvqdԾ��}�5���:��,"�1x�G	3jR�r�6	��/F����L=�f�>��y�$�bˎM�ه ����·��a�};�Ѕ�x
�5�$D�j�S���˫ұ�n�gq�h?[F[X�8�S�r�Z�zFV��1�0��Lp+L��k�]C�G��� w�h��ۗM�D��Rv���a>��jpPyHyp$�>빅3:8Y_�>i��5ҝA���6@�,�+�s2@i���U6 Q�6u��r]'�-��Պ�AJ8�����uq�$q��	��ᘧ5L�,^]j>�)9!v���a҅x��s�_h7����=�mRVw9��'�
[��qtI������퐡���w�%5g�q����c g�c�v�!����'�(�Ya�V�ē�s#�p��es�t5�y�����h�B���~��Vp�� !G!Jr��O�?Ctu$�_֣��p�{b �Da �K�I8�Y;s�l���=�������ȝK ��|��b�r��s�ѳ��O|^�5��n��@P5�?K��Vf����W���� �G�g�e˲Z<�!�"��lL�)걢�Z,aj��0�ܳ怀
�J�˿�C��������v(�_��2�%uuH]�_�r�A������zY
��R}����W��E�PCeQ2-��� ,H/�/НV6*��G��c�������ť�!��i۬����χ{e�\�V#������*g��P_������<m�/��{�#y1�X�8셢��M�����	��PjB�0�p묳���t�	��S�ܑ�svS����/��퐝6��Dr#yd�Ĩ2�)�����bT-�~&K�{�������� =��m���y��^J���^�J�"��J�>�8�4"���S��H���HDRx������kߺ��B3?��P���]t�LA�����I��&�g0{-�#��Oh�si����Pٷ��9w�Lu �s�0&��B�~O"�6)M�$�T������Ξ�����J"�\J$���^):���	A,{��EƇqҟ��@��hY�ȨWt�-#���Z]}�:�L7B�P�l,�d
�@-�S���!=8�?��U�����1�0�-l'Q!�;fJr��y���ð�Fp�F:��� ��{��S��i���8�6T��c�1v��&�};�Z�+ݾ���SZ�q���Gm�i�Sr*�mj���pm^�ǵl�PAt��ga�i`�%/��D�a�]�?�C7A=�o�,��B$�vp�Պ���EƐ_oѾN#H���Ƈ���"�/���y�o�2@��`"�˷�+�*�e��>��ᗟQ�]�̡~�R����p+�K��C��_1����`65��uQJN��u��\Hb��ܮ�M�KH��q��Ŭ0�kc��l*D��#�b/�䧁M�8^J7��$�iU�H���4��q��"ߍ7�����u��>���5r�5��P��<�����~�7Vt���
Ħځ�p�u�^�!�Q�ŽU7�@��#%�g���}�߭S���>��F�	h-U�8$ò+�i���3�7M�9LK�i�{c��23���w�����j�ͮ=�i
!�f�)�|����!���;ؖݡ4r��� ���Mhxw��w���R���!˄�Qe:y}h��U��o����:%ŭ����6)Xau�7�%W�w�_���,�k��Wo (�f�U�b7ws���o�q]���i�����|��E曞���
i�ޅY��@��5��H��l0���`�O�=2}�W�ARm�M�N��jS��,�Q�3�>�8���߀�n��s��]o>�a$ybnA�Ȭ�ԁD��[��1.�;��a\D����[�.D��έ��(�}����#�%�y�I���s)�f�cǪ�bnC& �n��O� �.�?>,��~7m���	�����,�X��@��$��;@v�詁	�c��0���[�uD�#��T�^\�-���es��W0�Z������Т���i*G<)J;Wi�v�rB#���}ۏ�H��(h�zI������ Xx в��^h4��p�	�����R�w�b<9�0р�i*��i��Y�[����֡F�����ge3!DG2�D��9��۷�n��V�Ԥ�k�n?�ЁJ@����S\[��[7��9��_�WY팈���k��]���Q)O����|���?M7�k3�N�3O�M�-��p����Z)�'��YQޤ�6-�ԯ��H�Ƈs�]�^,���_�쓭~+��E�}v���HKә�/����
�K͛Fe� �m�d���$��ǧ��E)5��8��J�=�ʦ2��(F���i��}d��~�~�`r�8���+|�� ��.4�������<le�(��C����2�蛮�O>d�5����c疼��K�dUo�Q7P�n����̓�Nʩ����Y�*i=�4b�*��� �v�3E�3qO��J����s+�F��[��ߧb=@�
}�gў��t3q6oO�exw�JjU�zPI,b⢉m���i�<�Fޙ�@�XsuÆ��Q횶��o�@��w�,}��T�z�24��A��� a��B$���AB8T���ND�-8�t����=���E%����\�5�yGGU��!�m̊����T��I�R�IY��&7���T�=O�d�\B� #+���c)	����Ox<�`$D
>/B����=�E4��H�g�y�A4F���|䴵H$��������K�D̆*Q����?n0�.�b�E��;s���-�W=ò;KE���ȧ882aMI�/����^�Jz��W�1j�U��_��f0��Mpy<)����~i�$Bh�'�5��xsK�ᅁQ듧��;�ɿ�96��qoy�$>;o�z�ZQKʫ%���{+�O`���!�����H���GPoS��<�0N���6M���/	����c�O=ęҥ�6\�O���C��J�u8Z|6B���+\��� Ct	�%� �O�ܯPx��(���+�%=ib�QQO���pB�
o��T3�O+r�k6v	�s|U\:I
���)��4��T4�0�!#�ٷ8U|O�*A�hB,{�)\�������i�^���B#J�Ic�;���G���o���(V�:�i���WG�̮�HGy@S���1��gl��98{,{>S�����l����-|��&���3�I� F�ആ�%T�I�Iq��Z���1�vևD7�V�M|'��N���l�x&�ri�Δ�7�+�<Ȼ�\Jp���`1[����_��c��WX>�b��rLmD:��YERaߐԊ)(��ϸ6�E_Z��1����DH;�x�
Yt�'B�~�%���U��{Չ���x$��iq�a��t�A|��R�[$�@�����ww-�,�d���������9U�w��ͧCj"���o.��ز����e̝>ػڷ�&��ro��,Z:��_�]����0���%�6Ml����'nGMڐ!�N��cw#�璳��I�?��xd#�����W�f�֔1ܽa&�������51�UfS�m�+��+o�F����q�ߞ1�� ��H�J>�ݍ�8B�����~���2�ph�=`�'����W�7��ѕ�A{���C}C�� �ђ�����x�~Ƣ4/��� J��B\�6�^v�������U2uq�U�� �).t�W��J�}��ξ��էvEQ� &d�,u��l,�h譗z<�-^��}[��◿%`���#4�Ϥꍌ��I;˗O1�lQ�`�N}��A��7��)��T�4���#l
H=��U?;�5�A��+@XS�e���j�-�%��6,?ίS��yK�����aw &��Q��&	�n0��!�>�����y���-���!l����|$FHZ����o|v҂i��
@g�	�7����4�ZN]�p������ʙ�ݩ��]1�;J�Ʋ�3���J�v'I�A��ٝӥ�\�e`�	�c=�q����伣� ����w/�Ε����=��<_&���G�<�0�T)�,�J���֦�,�_��4KC=/Җ)sױ�wo�_��~4suso���;���,�q��7W�y���/��d� �L:�D�C!"���=������ِ�:��m�2%Y��},��_4���I��%�pV�Z�����%p�Z�Q^����	n	���������X7#��s��)���<�!���<��^�(}��rO#�V���deL!�`P�T�(G�*��N�ȃ8��:;�"��1�(�uw��4�aBBd��y�7�r�hλ0�_k!+��8���Ji���
8*L�0��ލ���,]j�#��Mg(D�-�%Ь"zY'�qh����r��	�}a'$��J��PFS�A�@m�߃ח�D�#^h�)�&���"$@�o�����	��t�];����v����E�.st�R��]D�r��=�+u]�y}����I>�K���.Jm� ʃ!T�qs�{z�۩�&s�I���X��;V̱TUD�|M�����X=���R3v�Ը��m��IJV���k }��B�-��hʾ����v�"�#EO
����-h��߻{o5���ƊO��ڴ�\�<�sC�%��<�����ʄ�<@���8���v.���8���>�[�40����D��o�f������CZ�)�ʩ��Asq�ʳbLP�b���ۇ��N�^ �M�9���M7%Hh(�:���������g����Q��è�5�B|�e����Po-5�P�1�p&tqߐ9���Vj�[AX�W����w!��$P����S+"��h�*����OA��J�V�<��=3(�c��m�������b����r��K����?�� �{�C!�_]��<�KƑ�~R�Uy!+
�[��cRc\0�k�\���{�u�G_C&���1s)԰���6��O�ަ�c�!r�r�����wCW���k�����jvC�Y�.jcI0
��vR�+!w}�,V���|�����7L"P���4�md;>@C�QV�zJ7�OE�o\b�����u�����I7<��	��8��~�����D�zݫ�0k@ѯ�`<�8@�c�ⷙ��:�=#�1��ۃ���˂�z��ҙ&���g��z�?�1^Htÿ*�Zv���u�2O��C��b�Lkј��	]m� B��@"&��1��IF�C?=��?m�����B��ŷ"9A'�*�H���d������H�6�z���B=�����l̒��GF�/"��hϸ��If�T�U��u�Ki�$9���ԓt`���%¦i��W/����X�,��_
$TM3�ɑ�o������R)�ø+T�x#��m�h� ����Dې�*�AV>gQ�U�M���9�0/�? �L�a�ɽ�~��7����՚D9Z�Sj�i���y�����	���A!�C�׸�qn�a�`�0��_E���P=y�l�,����0W�	��6h5��D5=��s����_��z�>�5w{�
�>��J���L�s�S��Х�4X�+΁���B��񢳾u��P+mH>�rm7�yN�=�D��8�{ �b%�蠟���᭟#4���%���`Ȏ%�7Iu��P�W�諀�-�� ��B�T�@3ݵ���S���h�<�\�Exa5Ȭ�'WT�7���
#�d~pK�.�<D��8T��k��[�]F$ĕ#�&���܁\�z�~B��Dz_�V#��'E����]/� t�1]9���O��w�I�����+�d�dR���,�Y'nd4꣚ȉ��߁�Z���Khr"�S�.�+�l��?=���75s�Z��Q����9�\*�V/��ɋ_FS�b��*��7�'�������aR�"�������r�~^ö'9
��C�B)�V����8P�Ȧj�'�}d.����y<�4��3�X��l��ؤ�Qm����#����ףԲuMvB�n��[�B#f��P�Kx
�:�IJH�����(�S�x�C_g)!�|���M"�ϝi�q��:�Y��Si�-1��L?Jf� E agZ��\�A7��_sX>y9���T��3�9�}�~��i���^�4�����sRQ�vq�'b���G��?����3�J�D��-���x�[��~Eɫ{��n)d]wb�~�+G*�!��$3�Z�W<��m7��:��h�2�/(��yky�8\�Ǧ��#Q@���T�Q����w����V-V��s�6�EH��t�A� r����{;j�1T
j����޵�g۝>�O_��C.i�88),�]�����Y���,%�J�F��)u����Gd�iH��-�V�U/!8�#(Dw�l��\������C��.%��@���l��k$Tf�C"�����;� ��3�TG��1��I4^8����j�$�q�%�iG���§k�a$B;'䎏5�#_�X�`���������{�2�oYC~
�m@E�����oe��`��`��<���Gji=���ޣ� vSf��o�=:ԲB��e��NA��ݘ_L~�+C�K�XfS��鋷 F�I~e�~/��g7]نo�ٷ����h��c��0����L��=�#r/zýE#KLlo�Ƌ��hҌ��9�ם~m&��X
v��?��]�N��dW7c��D�YU�2�S���e���|���l��s%M���61�v��C��+~����%3�}"�J[����	ޚ��+rrܲ�'kZ[+a���P��9 ��P~꒡A"�W>�P�_w�G�^��4��0>�p3�3�ǿ(��C�Hxx�S�������xf���]�Bg�Fa��Yþ.Y��4�%?Z�F|�f�U7��i��8��ɵ��ٮ�Gfx
�t����I�
�q{liJ�k���Rc�▿/*�u����/�j ����ec�����0����n���� #��kC�T��z33@ 3#Q�X�dv����(�%��xb�ɣ{��9w��u=)�fՁ���Ch^ @Db�^�ɛ�b�2 g��G��_�ġ��sU(�f�	0�pK_h�� '���h5ˋ�\r�^D���_�c�͞�#j�J��zA@��)���5�W�_�����,F����n,Im�˲���
���{m���1�L*�k��*��*�/*h��tTr�i�i�m6�|��=߶;6W	F���9af`�[`�Շ���Z�sf��j���jX�QEp*���,w�&,��p;ݠ�kJy�k8"��n��O�DS��"��)VY�J�9�ά�$'V03)�4Ιm�:j�ԭ�W��P��F��C�[E��8_����G�H���`iSߐ}����V�q��}�>�A��8Ev�J�����؎4o��ɭ�".^:SX������3�z*�\�6���E���BoGl5ĽjU��$��+�g��z���407f���=���3E�ۄ�0�Wv�ٯ���B�=Cz�d� U�َ��	0�����.��e��b�T�B��e�n�&4(0�vͺ�p� ��\Uxĥm��*��������/����
^���;�RF��2�d5��*�� BJ�
�b�9(�fs���yP	4����7��4:0��i�Gu��60�&2+�Ø�D��UAf8��8���N��u���qB�����'����"��Mֆ�O`en�*����QP���1��ǩ*����o�Q��ҩ�B��@�$�c�v��h����)�[�������}��!�,:��#��xTH5��|7�h�V�Ej�>$��%.��~c�y�/�����%�?ۗ_���t��`� y�88@��"������9�)�����RZ��	�o�IZ�4�/�K����:�����\u�#
F�,e�j�S�X�QC��p?���Qaj�~�Q�s^^�߽yT��K��tfag|����c�O�Al{(}"�M�P���/��.���+��^���ӎH���0�o�Y���ԙ���UGd�en����<3,Ů0|�}��e3Yq�օ������;�W�;`|�4�H�M]#���&8�Ϡ�b�!��Hi�C�?W2�pea�)�A�O�V*F�xi����=8oX�v;�O=g��kFtaE	�/�]���X0b�f�2�1v/��XT�����909�g��vQ �F\��(X�Wa�F��@�~!)���Z�ZT���*�S����G#��3�'�P����>��K�7r�2�%��,�\a�67�c��XRһCr�BY��^�JU�_����
-�$
h9��G��I� ��s��sS�̘,Jm��o��w6sNy�Zz�˾�n�lS\?Pc�����Nz��.	D�J�%�W��?�S��X�0���o|q����� =�~ɱoӟ(��1�/VF��e:�d�_s]�L���@g����T�U`�ae��:������ǡQ���$6�H��B�/��؁͇;��Fg�Z*ezHU)��#º�F	�c��w��E�ɯ'���:%ING�Wv_i�!@Ԟ��$NK~ndOl�%I�*������>SJ���l�ق�� |�,ָ�Pu�j���їĊ�@U'��p�s�^*3)ɵ�5��?�>���x	��c�9�+
.�Ϝo�[K? a�В�R��Il��K�d�8?��#h��
�}���l�<4&� #֣�yW?�
�f>  �������A�W�H!Ɖ�ŉ��G t�|���1��3��r7�����ȝ�R��I��%���o�X8��3�E(�~�%X���RhP7�vj�{�ݯ���4z�����Tm�65���k3�����e+���\s�})�tR�ΐ?Ŭe�����n����ž�U��\�D�-�c�]ʑv�a^^�)#�m��H���~؋��DI�C��).���!t�+G\��#��+1��x`#�-,e�૙�WZ:��G�)�r��t*�K�Q�l֏yʉ����A�`˳���WQ��wC�V]'��NRsmn��	p%�}1V����`��V��r͖��[cPB`�oS���X����3��X�E��z����~,��3O�lP%��?��Q���i�̄D��h���^��U_>���tMTR D7�����=�!���*�*G�]J��>p�\�K��1\�!�e�	��y�l=&�Nj$�LD��Bl�J�ɴ��	�8���z^~\�CA�+z\��N�b�z.d)�A)~1d��t�Y�
�|�s��B�-*��r2>P������ҭ��3��&�M�ו��̆�j2�C9M�W֪��c�At�ɪA��?�Ý�)O�[�5<�՟�p|
c8�1�<{-�e?{_�o0��'8�
�}���dbB�P��V0Ϡ:�r�=$?`w| ��yH���ӵ��FC<�.\�p�fڹ� ���b��FF� ��T46T���Y�O ~�*���C��Q�S����0H���d\��Ќ��j��Z�����+���"�w�(�I��g����wl�q�[��A!8"����/
�E�1v�3�#��j�
�,��/�5�W�:�jU��{�G��/'�L���B'_��� 3ZT8��=�fu��\Z��~�>�9mL���m.\��9����br�`q��u�����Cx�IĽ����t�%���6��F� ��wTH��uN�����X k��Tٚ�x�rd"�^ʷU
��g�^�����wHff�bD4U3vس���Ǔ5v�w�/�9��S�-��K;���R�N��2�\���j��H�3�ɣ^�z�� 2��5Pcv�t����K�q�={�fZq��ӫ]����# ��?XOtH�D��P_�޳����^����GX����!L˔�3VV�X���.1<��os߲.dL�W�I�F��;Yf�k����h�8�YD��My-eR�>���}��}T����#T����ѿ}����dŎ ��3ߺ��P�P"}LQu������4l
+9s~���	��_�
h����������R�kX,���L-#q��l7��/ki�O-���=#K�#ڞ�9A�aʸ��wH#�M���F�mrޟ7���qd,(�Ȼ[�̃���\i��i��a�I<���;�FY�ȼ�>m:���h>�����z�
�P�ɻ��t�;��2��a�?vmy�2�/�0��P}	����5;�:j�(�����Wt">X=
��P֕
�Ώa��:L��W �9���yk��C��E!������J�"ߜ��B�ϔFK�9N0Q3�J���k2�#V�e��a�?��z_��ds��5�k����]<D!����ZU��h�\宵#��钍��!�d-l�Y��wT����'U���H�2!�C=o3�t���X��_�0����x����56��y��E��.�C��Y,�>���Q�t�4{�O�6#��n��>&����)I�vW{�sf1��j�=gm����0cE��c�<��PX�X!A��H >�En��%=��U��0��Y��#p���� 8p�@���+�aR&6�bˊP���?�l&s0i�~e��ʮa��'��M�e%�L���Ο����ݜ~�e��1���qj*&k`H%L?)b"�� �Q�JrG����;�G4��7�/�{���f�(�gt�b7�m�6L[K�;f��W�ba���}�b���{3HN>�q8����rh>6����x���k!�ImԞ�I�� =4�iF��Ԯ�"ty����P<�-YA��_El/�8���x���*�Y��:��%p�����i�p�/X[|��KFw��<�n�����7�X�
�`e��Sn�e�Wp�$(Sk��1��_�91|<mt/���$sL @�	t���"ys<�lC�2��~��^ԲHg�AO��S,��f9��Wu'|7&����cYX�[�.n��}FW�<�>�~�!fR mw�K�_�t�}��������`�k��b.����Hq$�&��//&b��(;K͸Hˇ���.�&Qfn�"`s'+\&K>��&��j���cO1Ɠ}*UȚ�嘻|e)I���{q�BX����y�Tʲ��~Gtv�=�-SxDk�i�1�좭ļA0���_�¤ ]�i�*�g��>�Pޡ�3��D��1�-�<#!fSIj���bWfM��03(����˿���'?L�*F	�5���C�ي��3ܤaʆw8�����j�G�5j��6y�����Rؕ��h�e�w�j��g��/9!#u��u.�b:^z�q�?� ���)]��'ϋ�C�U���2Z���Ͱ����&�"(&T`n��;����_�;?�K�_���eE&�wa;b���d��y�[`�Ga;*�z�9 j���gqq6ē�&�$@?�k��4b���X���O����%���b�R����?��&m���i���BN�M:x> 
~����UO�¦�@4�B'�Q'�6y�zjC�ke�cwJ�qP�݅Q1u\_v����<�~}�H��L�.�����Q�_��f���h�Ӥ`h�F�Y�	G ��*�Ne$gF�Q5��p^���m����A�q{��, ����I/��B&��1�T�i̱d�׳b@�:��/l�V9�0;�*-���{W�X2���e$7E��S�қGo�~c�-n�O�W��,Sx��l<�k�Ф��X=���#�4���"&F/I�8�i��;���L������
�k$�������/d�y��D_�m��`qFO��$[�	t��/���<_�D.*w�)e���	�ֳ�
?�l%�6�&������-�d$G�g�b/T��Fٔm�� �j9���4=��C�G<_9�#!i�H�11���x�X���>,O��h��a�<�̝��t'^M���D���ECt�c���K>�N8���!�a�����>��|��})��5�՞�Ews\�U��M���b�
�7���޵�%�[��A&!�^�؊�b���mc��Y��a�'G$�<�U�Ԅ�?i�m��+LZ�,[gW,7�F���7xB���6�'�>�e��g�]�E�!SYAz������$ �K�&?k�^l�:h4���C�2�J7���+�5ע��)���kɾ(k S�w�6G_�i�O�
ߏ�c��>i@9j���Z�k�%�@w��56���\����(qRI�0��v9��x��Ð�x��l�W.�f��5�agk�n�f�@���J�p�zV-Y�z=���t�i̊%�1���T��2Jo� $�yu����r �ur�Q	{��/U�t9��5ON��o�^NW�;�ّ��+5��������k��w����	>|i֖p����mη�Ot������Wz����j��vF�d�ا]�
���)��|�l�h$/�����Y`դY����TqC,濮	�3dݸ�Nc�v':
w�L�^�$x�E��+:.�lx��-�?A���{g�Y�ө`�ʘW��5+]:��
�CD����8CU��ༀ/��:����CVQ��d�D3��}��dxڙ-g�ܲ�u2��?��|����1�H�yU_���%�8P�U�
΄ ���+�,2�^Jm)j�ʱkt�u��W7��H�̸�>r�qisO9�8�����,`�WIUB��=fX"�\���i�&�M���=�ml�ؐO��=�bF��O �NtLR��gD��^����w���[H�ܚC�~#6�+j؍Af�4xq����G�J>E���[�����O�/ӲDDR=�"gj0�O,����+��Ֆ����~�DZ���j����?1Sǫ��F�����^"���Yb�Y�5^�\1]�� �mu�9U٢k�w$Њ�o>s�0L��ڨO!���z�cP
��T+C%P�g��0�i��s�L��A4Dg9op���Q�܆�����[�k�g����1J%����o�X$�_B'y�C��|V���GnW��-)�jW7�<�T?y���.��-�k"(�2�\�,��������W�s1�f�5C/ݓC�4�F�o��鰶��^~@�	W��9��5�B��
�e�d�a��S��͊6V1I�S���T�͎�5Io6I�=Eh�&n}F�6�\��sM'�,��v�;����$�t'�Y7�����x���M�Nk`?������3��L�Cb43���F~���J\i��UʣP����ǝ�?�^=2�1C�s���n|��������Hk�T���ª8�ҟ�����Y�?�>���C7�����.��d7��Q���A�og��
�5��[(ʷ�8��wlzR!�8���w�@;��奜�V��Z�&~ _Vz4����^�gִ�z0��R\��_�H�h�8���꬘�2�S��#̪����J�K�u�dn��^�-AY�����Ð����>	Vȏm����ec-�|��y���0����N=�Oç����ɩ^ᩓ3��]����,W�-h�Pz�
�
(2}$�/��~bGN{���}�?�����!�Y؞Q��`����zB�X}l�#���M���鄭M��"��'�@�NA���ß�+�ض�?x<����Y-��RT�pt�F��Z_80dD>��O���B#��an�Ȟ�4��s(� qMò79B�l*vdIN��)9�5\��ړ\'S�
�YC�0�3�Ǩ�.�F*�!�L�!P�/)q�@L����8�t}k	ݳ��U;�C9��lT6>b�@�k�m�`J3_�aotI<�;�Mip<-<����h��ˡ��w�v"y��zC>r��&V����gl�J�����u(�2� �#��N�B���\D�Z��c�Թd%,����j�q�GO�"Aip�ѵ8*�ץ����o��k:�7�����0v�Q��8M��h��[��B>�X�[s��N�ji/�U��֩��� ,����F�o���2p|J�s+,sܸ6�^�c�'��M���<kmQC5>o�z{�QpTr�����|+\Ɋ�ol��N�;�Xǹ�K��~��Z��ny��ǆ	��MbZ���'��h��`�(87��W�����>,~b�k��4�9R�ǞB������:�:��YI�'�����讖I�� �)��[����R؁�b�?���;x��)�i]!�'�l1�^Z^4W�>���l4 ��yҚQt��ƪ�E���"�db�O�8�D$�I���op�����4h��
!���uӳ2�o1�?q_3v�OPw�FO���1�]�y��Q2���+����!#qЬ]��XA���0��0	$J������=C��Ir�D����K��nM�}�&�' ߑl��G����쬸���4��LSĨä���clY�5���>�g1�./��x�v�� &��, ��}����2�ۢ��Wv�B8��Yy�z�U�:DSm������&�',駫2$��% 	?��d�X�1�wKB����r�SIu���C;yL5�1N�	 E����1���v�N"��$G��M�B�>Y�T�6�h�ֺJ���E�S�����R4kY��>;�%���g��$��~����#����~���0�*C��L��[U�ir�qDw)!:_DQ1
�N�xs��bF�\��%:\�� =
��G��`����0q�˹x�ʩ�ϸY�!�[�z��6�$�b�3�p��F����O�%$�):��������La��>؍�$�v�k^�SC���������h$+���^�Q:������G�mj��7ɏ5�2hۣ@6�b�C�I�S�:�Z��&�C����'k�1���D���x~�Ϩ/ؙ��i �Z�YŠ�Y�tPՅ�y��R�A#0�t�+d�C��/���F�.6",:q�� ���\���m������@%�"�(�Q5�;3��\���a�ze��FE����_�iO���;\���1 &�Dv�r�Gn�tG�?���CDB�!T� ��cIf��(!׶�/��o�A�u�z�9�n\�Uw�n��Q*k��x9Ch�m�׋�}��(Mg�~���!��x)�!K�O��EY�&x��~�QF���o�+!����[��ϝ��X3�K�{��lO�B������|�Qܦ-�Q#4�!#&��3��oNfg	��V��A��0�Z>���b|��wI�ǡLz�����A`�-r��Ԭ�هb����3#�K���]!Wm,-����>Z�_Q�������R�?�������K�pqk5������1a�zݬPd|��k{��?�.x�'���2F� f�u��qv6���L�O9D�E��VQK�t��n����5��^�}�u��	�K�wk�И:$�l�X6�:�h �}���KC�w��Z/J�+J�%Ɲ��5[Sbl����ƿ�Y���r�z.cl-`���Y�j�z���s{�l4�AT|�s���T��)]9+�&@&��Z��
��R�BŪm�
��72
���M��Pڭ��:���4hk�I�U�#����6)���Y�&��B�m�E��o�U�S�&T�*FG��vF�L�YDI��.]�|�y*�i�jq	FB���y)��;Q��{Lc�gw�^���{F.6��D�X����RN�S�h�x�@!��t�TyLH�2�� d8�zA�΁!�[GR�R $>�,�[�zN��=Y,�ʸ^��[)hf�Cu����L3�ԉ��s���C�̌��j&p����m|�Q��
���)�[DS]�52l�1�1��2�����ϴ��pt�tl�@��X��+ U��EN�;%�����n坡�(��
�-8-�J�K����3=~�C
͞�Y�=������k���R()o�����Պ�^��$:�+���l����\�s3O�4M��xófս�a��3�Y4�E �!ghM���t���8x�鵙��dwc[�hm�e#��=_�<=8g�kb�b���]��Ƚ��)�W�o0��h�a_){e@�3k�0b3�L]��10{��H�_C��<:���֬ɶE�K,�����*�K�ܧ�:��$i����w�i�úN�����/ba�[͡,�c9>+��^r�%�`�0 ��68i��*}��dM!S���9W�-z�~؞dD�����{	 Uq���V�#�'cU%ۑY0U�3�H�O��z{�������n���{�>q BaN �0#9T�"�|�19ja[w����4����������G�FK����&��x F�T$��.�}wx�?̩��S�8)c����?:��gM���Y�qj��0m��X�;~��v��P�t���S!�qV�S�w�;\�G��	W��d[�ъ�6c������0s�G��J9�VA���1]�y�����{��s����
5#��$I��H�|���؁����4a@һW�Ȃ5��~t3����1%�~��>US��q��<x͆�M[���׃o�f	u�H�����-u���Z�f�� ��� ���u� Y�:��Z��wA���ُ<���D�b�a�����ѝ�RΠe,`�V()�(�+��@O�����+:�e
:&���BT�����"�e�eH�y��z��n���v�/�"�ow~G��K��@���!��n!���YY�RqwU؆K�\J�|��l��֑,f����$P@��RG?�ʚ���pN��e���)����N�8H�h&��M>d����M�8������ˏ5cz&Ln¾!���L�͂]#b��w�/��l ��blE�&��5k�聋�o�̅�K|r{v��� �wݔl��dp��e�t�U�xciu���9�c=V̌%r�7��[���w�l��?�����׮y}pi�t{�Qd�.�*��t2�|�-:)^�J�jAD���2ܶ@��~�zK��=�Ԃ�ITH�7r`.Te�k��=��#1�4B��A�g�� '�c�'�� ��?���2�렸
}M�o�Aĥ����\1\���K9��F4�]	,eq��쿊�:�{��s_�1�-ikO\7�8��? ��Bs�O�K6�L/u�Q����s�7W�V�����'�=�r��d��/4$�(G'ß�*1 ձ��4!��I���q�i����Gz�I�$�Kكa�א�p�v��.�*�'��B�{�'ϕ¿�Q��[J��B+ӳ�PMGF.d���/���<lu
�X����L�M�%x��AX�B��=����6�ĦYyI\�X>���7,�Ez	�e}���~�3)3т7s����C��  ��Y��(��?�B��v�ƛ[�j�ݾK��z8E��;��zS���a�����ԁ�R�C�l��ڃ:m���x��G:���ot��Ϧ4�sN�u�J���NIʘ���`�ڹ_j%8l`����F[\�*�-"�al�T�?_�h\���/(4�@w���C�Y��uQ+7��(O�b"'�q6zc�#����/�
շ~��m QVj[��2��HGo2�O0g �z�Z�&g�w���墶���#�&N�L�I���$�i]�n����워.
�d�6;bؼR��pB�b��Dv����QǠC�׿$�������a�Q�z��=ݡ)�b�f�5H{���I����� t����O�m	��W,Q�]�[U,�>q��"	���N�Q�&��٫6�@�p���F��Вx�y�=|w��zE����)��ʵU���X�P��&DC(C��PiW* ��'z��WU��Yj�m�A֓�,�B�vK�S� aR�MƐ"�E�9_��VƘ}��z("�ӹ��J�n?Q�/d�h+nSa��!bj�3�!���׳��&���fL�:��Ci��&�ҽ��y��(��<P*j��\J4��k�*	���h``��-26���y��u��B~H���j����H�ی��\._��#:�� R��my�J����S��|Q5�*yMU������W�Hj�Y�߽���:�3Ɖ���:x�i��R:V�������m1�,�(�`G��:|J��� ��p�~��;E�JÝѼ7��������J��'	'�f���@Sz�!���<72����������JC�+���Bg(����`Йeݞ���¿ًV���pl�T5�����7t<*��~��Ӹ�v���4R�T�)�>��97�<ɽז=�Fz��i�� 0�R��L��ڄ��p�>?�E�w�g��7�ʶ%�&dr4B�(�� 8��0��V��Ry���h:/�C?���8�В���N9"�����y� �@�[���f�A�a9��+�� |�i*Ж7���ę�;��ׄ\j	WS��l��m<��2&
���R��l7�=LX�47�#���N%�����U�mf�����8�l:vS�F�����p��2�f�F� �⢑���I;�y'����h�w{���Ө^!��9�ۇ>�>� �����7��|ޭ����n)�O�j'G�W�t��Xס�O	�I��^�����L�L�G���b��:P�=њ���^�t�'���G��&����\Bs|ΰ��R�UeP�����DR|hR	7 w���L�8t7e`X���w��NM]��hn.��9iP���|)����O�3�G���s���:SI9�O��+Ow�[N|�~�p�ƍI�����խ%�@���[c�z�3�47����V��bx����Sk�+�a­E���~��
�6�� �}�g��\�<d�ۢa�7k4���Xp�{�j��f?���.������+O�U��%��w��!�g-_��<;�JJC���\.��+T���v��ml=|�)N�5��`Q�f��P�wo�o�K�:��$�W�*����.�楷ђ9�[��u=A�>�k�d(�*���~��BP9>D�ݥ�#�ދ��Q*o�|�s�Q��w�/~��`�s5�����N �Ѝ=ִjg6�a��y�<�cd�zo��Ar��]�;,�_�����c ๒�+�=�$p�~��c�ܒ���6�Ďhj����l>8=o%�_v~B*��/�>����,������UZ�BL�3}��SV��痟�o��7����j��ǚ�������;4'$f9�lz>�hz����H� �\Vw��Ɗ���@:��]�L�f�Ye�@��gM��yfk/���k%�z�N%��/�"�6P���uJ�T������m5�����-0�S'��ڥ��\��K�ˎ/�׭L�Svk��m��#�� �b�z��v�b�/�k��TN���ǆp{81\%�}e�-j��ps_��{y���d�*IY�e^z���._>A`�d��k���9:�N����x�X�+OXÄ�g�!�����}U�^W��H������H�N������� �q<8�P����o���(J  D�k_�o&�[I)wܴ�"�)g�a�R9�kt�4�%�.�v��3dz��WfU`���˞j|��Hȴ1�ף5�:E�'�o���� "�K<�r�,}���^���إ
�1��L��"6�m5Ŷ&��rϥN�瘼�V!?}��T1. ��9 ?��$��r//j�q]i���$e|c�E?l�z� �� 5�O
�v@EV<)]&�B".����`x߂���b�h}��a�����-����8Ć~K�� Ǘ�������|�f������27
�߸N�T��GLMuӊ��9Ԥueԅu��%[W=�����;�F�{�����O�v5
�m[�Id�F�;ϣ%���,��=>��QL�B3�b��DXcu��J�Y��oCChEц"Zn����f�e��k��ax)�C)w�E)P�r�35�a(�1b#�zH4�Fl
�ZZ�U��Ӌ�5��H~?�v�o	��]�^���MH���׺�s婀��}�0�`]͏܃�+�k�`�]�y��<���p	�ӗ�w�jC ����Ÿo��9O����g�/d�\XM[ӫU@�;�GM�I��Ƈ�0���(*���T�t~��?�c�u�#����e�(*�q��֯�;�PO�SSv-N�i7ԯk7+O�Rأ�!I�E!P�\ͫ)O
v�'UՏ2� ���s�a
H�$DN82,��J�9�N���CI$����S��4l�4�^��R��ZP���u�@�5���¤�t�ske6�-'�R��hy+L��!�$��oF��VcpTa�K"H��(u��n����m(i��(^��~'�ÆB5���� �<嚓S����ˮ%;�{ S��t+��v�!D�\D�dc�zV��CV,Q�9����d�J��[����0_��o+2�P�sȍ�nH}�d�H��v��;.��kА�z!�T�bfT�e�jB)��#bũ�E%+��W͉
�VS��Q�������;���Sc�6՘��C�l�k���w���H▯�U��Z"U�6aU)%P���_�ԧ��	��% > �A�������va����d����r�!twގ�DV�������zx9Ý6�83���TdwG{�Ip�!?�������8�3�寈�p7�I�|rm[}������^�ח/]����>,B
�\4kx�� �שM�@��
<r�� ��� ��i�P��C�'��J�}��w	{��zYO����=\kU􄴗x|dR���� �ϳN�W�����f���o��g����@�W5��i~��W�����Vס��]	��}���v�GB3��еg�<<��6�pVO��˃�<�v�c�F��6o���\���m�������t��r���'N �FUcv�����
�b�7N䯓slKh<r��,D����K��6	e��W]x&�(�}�_�Ufg�-d��㩀E�qi�>ٶ�y�q�K�82R_[#��S���,������̿�(C�-Y�i����J3WY�/���i����b�j-"#d�|��Wӡ
\��v�[V1��'y�'[��c�	!e� Pr���?n��NI,�N��'X�����1�k+l���3����p�T�s�;��Q����TTʬ5w���>�oKse�X�5�[��Vf���{O���BpJ���68^McI=Ne|��c3!]���*�#�:I��:ܴ��$w}�hS��Na��6՟d�e0�V_��ہ<��g_��밞�7�I&d�&��㯪 �v .���`�gLu�h�q5�U�(�t*,D��j�1
����TG��;�-~$���x�����F�0�f�F2A�){5v#3��^Q
��|S[1��k�,���?<���E�]���;-��||1I��<�ZZ���7�L�<��������%s��,
g�|�@�U<�*tJ7v5�[0N{|�ܭ������?!�����:�-ۣ�����;���4"=�P5G�o���Ўn���.���T�>_���ޡ<\UW2�Y!��1<(h>eV�	�����vD���2ߨbϰр���#c���a{��,����T@+��EPd�Gk�)k�~�q�n�W���GkV߱���Rb9{~}d�����$����u?�[)?{�������v����<Wӥˎ쳯�s���MKT�Q�9Ǘ2>�:yھ-!�u��2#��R����y3����9vȐ�\%�Xe�h�y%z�����G�����1m���]�d�0m���V�6cB�[�請���j)���^�����;�ko���G(Q�Iv�ڟ�s��e/#���g��[�8x��[�KI(�C�� ��*��"�X����>���7����b(�±n|˰x!+G+�[u���=Y<Ȧш
H �����GC����I��U�k�H2RԚ�+t~ío�DZ�����2�2H�H�@�f�[$���Sm�J�l��>R���eoz�R!˳���T����w����ei�HB�wch�]8r��21	��gE�:g��ӧI��8Sc.��a�%�QHå���-i��<be8��I\̙��yq�����U�����Uc�5<eu�B��	6�0�7��hX�bS����P+rOy�/�	s�tD��`�1]�]q�FZ�1�9��1dO��nV�?Dޤ�Ča��z�An�P��"��#���9�P��W�!�M@U#D��w�x?��E>Q��3�e����ҫ��b�*������I���l�!�h��!��:Һ�p�-�WR�h��xC���\�<�"������γO;Y�K�����®�v���9zg��`2BɅD� ��>���b��t����n�K�d�[Y�lX�7*�>��c< 8pV0�9֎�Z�X�������������̛�z e���;����$ �DM���'��Y<G�FR���]0!�B1���]0U."��i��m7%���o�m��oɴ��%)�s�F_m��_c��:��t��;�sv	�u�*xH$�@}5a�7Eĺ�pH����Iq�M뻳P�1�CBA��IG�dir��j���ᗯ��
XD>��� �@xz���>���,A�̒=�YL���+ɗ��J�:�J-C�����z'��Z�Gi.�ڔ��A�J�2J��]�g��?{9�݋8��lۧ[�#�ӿ.�(�ʊT�$���Y��w�E�����t��>#j�	\I��T�o|O-���zRi��s�2�)<a��+R��ލ=��,�ɏ�j����G&�p�=(z�j��-��,�V�;�˻~�o���B�d�2�0�� ���op~��B�����s���O��(2R���[DN����6�!�ub�7Q bq�#x�Ѻ�;B���h�%8�t:{����E_:�4��\�X��	܆�qV2B�ʒ��Z�%=\2��`�����-��WW^�tԏr��3z����Sl�$��ο�:�e�� �<�U�r&Ϝ����/Q�V�ˑeT$p�BC���wrQ̶:��<rW�پ�����8{M�-{��p���.����č�k;,]4������)�du�E�b�����g`�a.��:_���-E��e�Y��:��*� ��jc�q�8��̀����#5�s����>��2�R����YBN������4�{[	�[�[��x�+j�ٹ@�g���%X�J���c�:����I;�ҡ���߃c���l��
�
n�k��Oi�夥��w�k��S5P��{��G��"`6tm^�.M���l�����L�4�S�ݰk��x��GF�ҜDX{�c���󳩦��f$�&t0���2�ع=E]_a�� �F�(n���mm͌��U��e��Yl
��p⒔ّ��B� ���X��-!�� ��q�,
:GÂ�褯�(��3�I��A��B����*��#�'4;��ux��.���M�yK�$��|��P�q�.�X'��X�Y��u
���͍�Ƶ�E�*22�l�z`��-�d�����9�*��{�p��i�@�
��!y���j��z��R�?�G�w�3fQ����uP�!��(�:6�	;��>:�$��������ɤ 0�ms���%��l��b�����^u%g�D�.�A1��@w��ez���C`�)��:Y����kAwU����}|�+!t�Ky��x~Qh>@�y
���K%��v��$�K١NG�n�]����*q`k������/�!�팤�B�P����v��G'��=�%��d���|3.�����X^���*�̀TpI�Y��Og*L!�NVG����g�,�&����Ŧ:�R���:�c�/��0g~�/��� ��ԡ[���Y�����rZo��4���B��s�,Wm�+S+�r�����4�a&k�6�z�,��.c�ݜ��.z�F�N	��&�����Cܛ;,�l�~������U%�	z�¿u�~�M�}��Vxe�U�Y���ޣ��)B-���?kc7Z�F�p4ti첉��97i<��#���I��
�P�Q�WL̦K��ڼ��$��g�����"|���pU�-P�\'�AO�b���T�J��5�5���-@Iro��G7f�,����[d��@a=�dg�c����B{�V�.^]�W"j�mH����
�2����J,��{��C�}�����K��z?����F�%��Y�сw�4˭?���g�2%�![�d	}�1�US}�mp�/z%Jd6�|Q�D�j�9��R[���\#w۸Gi8	\�Y|���� l���Pq���=���a���K9�ӆ�)��dS*��u�j�T�!�![j�)�]jN�:���cr43r��
e~�x.�C����:8����k��*�k�1�%�����w�����y'`:��.�4dy>�5���LA�J��U�V�3t�t KN��哭&����?�MQ�8���a�8�_�C�Ʒ~p �����`�<��N/���! �b�����2�1��XQ߲=�l��Z���G� 1��5�� ��@���߮�9�kCo���"�����m�Y-m2z�����l�D�^{�,�JڊB�㉧��qh�Ϥ�������wP��f$��@�n���_�k�o�z��s1�(Xՠ������K�P{��!H��5�;�N���y��iK!�O7z���] C�
Wa�����&R���{İ��C2)f�z�z�7 h�J��YDlPP�U�I��	b�ّ��ߡ2K���X�$��ۚ����m�LU]�%�27l ���P8)G˄�.'���x���Q,��9���|�F��_gls�����"��B
&����N�V{����������H��i����XUgr̜>��1���N�X췫r�ͦ��  ����
f���h��d�w��V����
W]z�yl4z��/��>�ġ�%�ÿS����ꟙ�T����;8Xţf&,t��'��-!�D�K��Bh<�)D�Ԩ�z�i!7im��q%4a�V�*��7p��� N�Է�'���m?��I�Uoy���"�ɞ��1���y�����Rs�e��Qr���ڼq�R_Gv��(� ?��җ�����N/�߭�{و8�xsK��� @ۆ8�$�Y��ɦ!���8��p{jTk��?��:v��I�y�B��`^Jr��N0�*��	��t��n����ݨBW�P�4�8ͅ�'=���:��C໊������n\F�ҭP���}lOi�K���AJc^�E*)W2�G���^5����I������=?J�j���1P-�����pF�΋r��23 q�
��j���-���¡A���et#i�RU���.m�٭� ��%)�����_;{Ӯ����V���b�/<?5�C?"=iH���rhe��GhР��7��X��~�k���Y�6s�c���!h��Hc�ޣY!B٫����� �����K� 	�Ƭ��ெz�[�!�����5��=�^�ru����Ʀ	-U2ua�a���9�k��$��t�p��z;�����>������dQ������[�u��&F~q.U�����0�} :?p*1�e����v���M�g���jjjQ����_��84�U��jt_a)[�Vv�34�v�|J���ln��6.��q׃+�`�J�w��LX�r��P��`�U�^�PM����Ch}����#��︗�L���(����La��F2˙?���)b���%VTtl����q��������v�pݜ�e��*�~4�K���aB��q�nO�fŹ��nn�lb�L��� �R]����n6U=2)9�P�B5%$��d����g.��Q/�ٵ���ha�L��^�4�b w�>�3g�d��g�̀��1��\ς�͙y�[g�$���W~��Zl���Kw���abR'�띪�����Ð�̱n�j^]�i,�1_j�����C�čqi�>�q��c�hٓ�~���󢆉�s(�X�m	��j�(!�̴�ʔ�je:b��Aw?���QB�{��\Q2���uP#��h��
�Q}���h��O���N�3��������2Z��
��t����i��Ip�ϓ�EL�p7�b��2��E���kҒ���c��p�v,���T �I����U���+e$��1��Kx�ܰ-znPb���4�0����9�3r���@q\Y?�}��o�T�/��&��~��SHK�f+��w��VP ޴��>�E��+���!��KVp�C�M2F��20`���I~I�V�^*�Mח�@�
ʨ_]\�@�z��"��*)O���`f��J1Yr�-�I5_�o�'Èr�!Ѽ�.�M�Y�Y��;�3k���.t�?��\T�B��Z�������#�w��}�nћfB�Y����P1�^g"�g�[UOJLDE$y��>.����}�~�L��	�GhΫ_<b�����o�G�7�`b����݋�,�]a.��]����C�B�Ϫ�F��T�ZS{�)������G&��q��3��t��A��u���Q�
u��ZI4ӖBǴ�����p��˿�lw��D�9�^z�K����\w�A����GQ'�w|�M�[��GbT��,�bF;���%�Px4L
��x���y���+u��.�2�_b����ۈ�$�9���n���/�։�KL�U�6rk��'ɕ+eK��?�@��Ae��C"���0�.��~���[����0��Y�9�E����H�+nV�s���@G&�^�r4΃?c��_���*���fZk	�I,I�G��_�|��5"��&�i��%�K�`���~���BCz<T�`��i���߬��u�g�a��W$��9m���0�h�k&;��B���Ёw��&�IUꄛ��H
<��#�$ �Y�>�� *#��5sa�!�<��$���g���
z��j
3��XDm����ѻ#A�rs�0��x��a6�A,h(%��T�tiKC�v\�+e.!��D��C+��蘐Ñy��%���?n��Oon��s����͌!�ߕ�g+sMM�5��&4����k �s��(�0W����yd�OՃ�9��j7�(rlDD���8c�x�����d�S�l����r��Ļ
�W��H����c�a���wW^�nQS%e,V3��	�7�%);����';^��������)/Ȁ�2��Yж2C�c�0�ח�d+G��Qk�GŤ �
�t'b�c��Fc�nٞ~j_�1���_��Q��S!_�m���J	>��w|Q��W�}	xW_B�G��=����2����:�$(#1A�c�
����o�!K�V0�6�(O��oe��$�jvNy�"���'�h�4G#5�KHS���Tc*" ���O���l�sfׁ`b�?����Vi
FhҎ*ϩ��
����"s�]H2�^xT21W1�@��lZ:~Z��ۋ�"�}d��L�Rr��xjG^��!l =V���ɹ �A��2��pa'�Ey�ᦩ2�CVܾ�n�W�=i4t�#�>-��?��T��Ї8��L��]��!O���T��#|��"dUZN��Dh8�{}A�/��;HQ��d
dy���f��5�!��(�x�z��k��P�3,�����1�Ȑ�Դ\gLr�d���"�QA�� ���=��!<����	Ls�r�!y��y�m�+@P75��lA{��ɔ~�t�q�3e���j�h�o>U��Ր��j�ۘ6u������� ��K1�ح�f���_�6н��
_!n��¾v*�֤���TN�����l�ΰ�H�$�d�X���-Sf�D���P�{�{�D�3�9�+�x-܍��57~vX	����n�"c>��_p��u@!��:� �U(X8?K�q��d��T)ܷh�m$S�A��T�t�:�
4 [ ��J2�{Cd-{\���eW���Ia.��C��Q�:��6o��<]��@�{��Aag\(Dg��_��Q�9��5��錎&�aD]�ť}�?M���.��\|�.��<�
\	�����I~΁"� ���dPc�q��t��T#Q�ةufʵ~3c�z�&$9���tB~�E�3�y��~C{A�1r���_�Tq������ݱ��?M;F�)�Iyh�k�E�i�-?��ֈ�v�:�-!��Q�����2�#��� �S��ڎ��7��S[KFz3"RGy�n���P޿$$�푌U�И����k	l��u�$��,8�(���x��dSg��S7O�5��]�H(R���մ��7�|���`3u�cv)�Uri`���1��Z��o�K���R�K4�&��dp}q��v�\����*�-�(�#���bgQ�(�� +��O<�m_�#��5�a�
���/+�1�7<j�i*��g�����v;`�ģr�ɱ{�rM��iVk�}��Nh��y���:��gg'Ȳ*���0\�qM��f9�?~���؜s��H%ר�%E������QS���j�@Į�^�zd�-4��:�Jbl6���-b�Â�E���5Ф��D���2zV�� �J| p�0�K�_