��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�\�� ���K�O�{��׮���^�ן��A�ߙc\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\�]���џ�_�v%�]��4�:j�l�,9��I{��8�H4%�}|>���ؤ����2Ee�Y�R2
�I.��k��[/�!�`�(i3ئ�!G�?|lw��JF#�+�o���B!�`�(i3!�`�(i30�mv�a[�y!�3�'��sȸ�"rRQ@w�ӏ{2�����Vc2�����Vc?�٩o
Ή[Ed�+��J�+�2�����Vc!��.���jsȸ�"rRJ�a$�Y "+��<k�K��;`|/2�����Vc2�����VcN�RPLo�i��ԇl2�����Vc�aW���n����y��4��ʮ�:I��� %M��z'7!�	?�">�
Jf��t�c�.[K��m��ĭ]�	��B�j��h��UH&��?�ї��#)kP���{<��ha��׫��Dx�A�c���>��k3�ݑ�����Ic�"K$y"�hA	� ^��y�C���"���87ۺ�Y;����4��Y�jή-��8�#���@�v�>H@����A+B�e�u�阻u}�����!Q�a��*��&�Bz�$���ş@�t�k��V�W�a�{Z��h� c��(�U���% 9�6�'Mcö]mҢ�Y=�FD��}��b.3O�C�L���u��Z���a�\�nyU�-�Y@��#)kP����:p#e�C �@nk���0�r ��s���̴�uS4My$y}�'^'��|I%�&זds£����&����q�HS|6h.:;��<�..�4��N<��;���u��w)�S-!������~篟|�T��/%i���6�ЛL�џ�_�v%䆎�[�2N�8�#��q�)R������}Z�
d~g+#���e��k�8���҆�|n��I�� �U!Z���������ѕ�������ֈ:Y�x���' ����l��m�!=�y����h�}�Zn�h�+��>iG�ɹ�6wx���Sd,�ϱ�ϖe��!h~S܄=S��r��~��e������k�8���҆�|n��5�ɻ��Ͽ��b~�wf��Df����C���;���΅iG��w�վ~N���m�!=�y����h�}�~߈#���0�.�	�Z�@�@ OK.B����Ҩ�j�E���H�ٳ,�M(F�N��d�>�l;��r�O��C��0��?,*���S��I����)h�D��'����!�zg�Z�$�R�7��P4<�`�H�0�Is���H&�dcY��RL�a)�ƞ��U<��I��8�J59��Y<S#-*�)!�zg�Z�$H�2��p���:n##���Ψ�	�ǳ�V)WϷO��(a[�d����]	i}���~LɈW��^&�K9���v���y��֥2���~"VL�r��=1.	+��(F����"�����dhV��%C_L����c�.[K��mN,����0j Oag�?�4�ʗ
� �AH�T�t��3��e��ME
��偀6�=$��-�P\~KP��:�h|�m���rR|ӌ
r�����]B@�v��8b�m�!=�y����h�}Y��݅ 0�A�X"zB�j�ǒ��Sd,�ϱ�L���Qep��p�R��$���wT��xݣL��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ����±�h���v'gn�]o��in�m��+�<4��ˌ�ň��h���T�%�/ң��Z����qM��D�J����S��������Ǜ�>�xj7�ܥ��2��O�����ϊ���f��8���� +��u*K6HT�����Np�S��<#l=���E����F�'n�^0o��~+�ݗ���3^�����n����\�v�e�g����\Y�4Eb��Y{�o��eŭR±���]SBÀcۄT�٥��T����kF����K�ca�?��J��Z\�'n�^0oM�D�;��-e>����C8�����M�g����!�`�(i3��|g�Y�'���Xw��������lԇ�-{�Y%T��BPe.��xu	�>��l%i�-ʲ��U�4�E����F��j���0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6����^���m���>!�`�(i3c��Et��q���U��>�w�Y�#� ����������5	���]���>����C��"��K��~f�[c��Et��q���U���
��I��N�Cٺ�������5	���]���>����C�/$�ߺ��]�P���Qi��(�
t�ژq���U�[��N�������l�
H�w���]���>����C�pॻ}��!�`�(i3c��Et�Y�{'%s��.|Z���ǚr��y�_��wBW��8���/�y����\mע������Y%T��BPe.��xu	�>��l%i�-�Wv�4�1�>��Z{����|g�Y�'���Xw�j�7��a(􆿳����^��/Z�o��>��Z{�Ǖ�(�
t��Y�{'%s�ui�铨g��U-�e�,���6+����3rn��yn_Fu��TD��ό���.�>�Q�c6�`S��|���Yl���#�]�!����M[��Ǣļ$����"�,�>E���TD��ό���.�>�Q�c6곍�ٜ�]Yl���#�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳����^��2�0���Q�#<4^���(�
t��Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9���6�e�:r�"J��M+7EEN�p!!v*!����a0��\�ټ�]�����q���:�0a�0��+3ǆ/������}	���w��Ot+�z��7G#+��\w��0]�m��
��1���&���]2�y�Z鎬���������o�	�*ZV)�J����67G#+�Ǘ0z�cUL|�]���?.�9$[{^7��y%%\�HP@�a�~�7���� ��JL�N{a�9Ow�Y��k��ı����V���}���s+����Q�Q&��������R(��z�j�)�q��1�:�Ω�s8�R�	�}�����ֶ�#3�Ba�b�Z��dÂ���dט�w��^���֮�LV����,JHn��z��p�Sg�3��ʹ�q�T�c�$�����2T�9�{uﱶ���_��a�\JS�Db����}�
�?�|� ���ܲ��+�J�����yg#��b!��u፠�w�`L�v�N�i����:��|}�
�?�pॻ}���'�gCm;�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳���2����.�t������ֹ ��ˎ��U�g�q���U��@����gG9�'��A+OV��#��6�d�٣��v_���Zo��`c�N��nrm؊(�h}Nw���}p$_~R_kV\�헌�]�!��11<�InN4�%;ך��C�:�S��0: ��q��MR�ۘY�{'%sAX���	q�KS���K����)��T�\ ��i3�|)sՀ��R�A0^L�H�߳Mkзq8�Ј'���Xw���,D�C�:�S����"c%�B7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���{.[��(��Y�b�΀�e��Ek�Z鎬����t��LJ��{�� ��8D�N������Q]� _�rs�i���`�M�	=̞��>����� +'������݃�Q[R�7}ϼ 8�������qJt� n���]�!����w�Հ�	�-�_Y��r-�T��v�z��]'���Xw�j�7���S�ڬ��M���q�tt�g��U-�e,%�0g�����9וP�;6�2�)r����'���XwI����"�d���m�0: ��q�"�k� ��Y�{'%sAX���	q�KS���K����)��T�\ ��i3�|)sՀO'�[m%#n���R�7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���z���Q����by��Fзq8�Ј'���Xw�h\K�5~�Wv�A��2���HF3}�
�?�/$�ߺ��]y�ei��nZ鎬������_�,�;�7���c�eK�	�$V�7s�9���o�jƓ�[b!��u�lv0�9l7s�9���o�jƓ�[b!��u፵�3i���Y�
��<�±�sR�{F�(R�?��f�Z��Δ9SF��.S����%�#�ڊ<?@x�����(�F�ܓH�;G+�ه�ݮ{�30�����ʍ��зq8�Ј'���Xw���,D�
�eM�6��`�B7d��n`5�fK�\w��0]b!��u�7�UyR�j�=l���]�!��	Ǹ�y85�����3�|#9���b!��u�s�Uo������zL�O�]�!����w�Հ��I��JnSl{�]&"(���+�J���q���U��@����gG5m�E��P�|�Ȝ��7s�9���o>��l%i�-��s=q�SbK����D�7���`Z鎬������_�,�����?�!�`�(i3%Ah�%4
>*"v%)��2��������� +_�XF�%�/kѶ���� ��Y�����E����F�'n�^0o**�ХM
�nGZ��JP��8\�S�.}�
�?�Y*�Ld�=�������d�٣���N N�S�qg2�K?\|iQP@�I	зq8�Ј'���Xw���,D���S�!�`�(i3�n`5�fK���Qi��+�`�������H���,>$�p�{�㘽2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��$O�a��Q�ڃ�)oY��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcZ��O��<�"��~Ǣ�)�s�ި�/$�ߺ��]�P���Qi����$~@퍜��Y�ؼQn!���Cs�9�+��N�5)��Z^S�QQ5��:ux����7��f:���x��
���Va�%��jq��/�a?�Ҟ��wɟs��A��e�����m�(1���&�����wɟs��Y�b�ν�r�� ��*ZV)�J�z0=�_���T1�8K��}!�#�b�Zj�|���ghR�P¢	�B�d�ZtgQ�9OZ��Q>ml�,"�x|ٲ��I����~u�g
�t����Zj�|���:�rQRт¢	�B�d����ψ/�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-�����*��=@rTnG��Q���;�Ӏ����QS��N��̉���G�+J��d�,1�!� ���үA,�&c����Q�nT ��{g�z�È�/&����� B�&"3݇F1�k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������7�,��n6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G7�wtMMP�~�9!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�Y������-JF����c����F��O�\E�W��4b-Ukc��R*SƇ���P_�2î��
�Ƈx ~����Z|
�Xy|�W�8�QeQ���{�`b+���Ãlv0�9lf�?ǉ�=!�`�(i3.5o�fa������������W��0M�Ŷ�z~�_m��y�i+����v�м�/!�`�(i3!�`�(i3�7uw��8�#4�?�G�{�`���φ��<�6�=�Y��q�$%��W����' �Ϟ)��K������f9�&U�)j�S���ܚ��@��f�\%`>��s�;�jmT�#�0M�Ŷ�Eʨ�`N/��n��<f�`u0�F��a�Va�ir :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3����-Jg8�iT��*���a���$f��_Ub����pT����d#�����"k�jCH�d*��=����h��LAи�����l���KyX�X:�^ao�_"e��� *�7s5kL�G��Hb6��l��� �M/*�3��7ݽ��x(�i��/R�ݚ�Н��k��M�� ��F�����@�9��n�7�Y���_j�����9�x�\M�ݚ�Н�;�V&S�b�4���n��Fr��jL��[�)�jMOBn��akz�
1���;��x����2�K��n@�Xy|�W1F#�֞q�$g�ޖ4�3❲{Dx�%�!t)�!�`�(i3���D4FF��&l�--|iQP@�I	��x���^�Q:��Tא �k/�ݚ�Н�!�`�(i3T ��(՛MSc����h��N�M�uz�M�Ӄ%�K��^/p#��I2�8��[�@����`����ݚ�Н�!�`�(i3�����zO^��;M7�`(>��Gƻ�������s �Ա�[���}��M�?L}�7�R��3��
�M����d��-��! ,IİB���_�ي5H�u���������Y��
�I�8����q �H�%��ZtV1{,�m���OG����ֺq٫[���%��Yڲ���g�Hמ]�NW�yߵc�Z*�NvM���Tf��tk�n3<�U[i�G5�
�&��zq��"�����¬�/���Sm[o�y'��BS�͓O�t$��Ŀ�R��(�>�N!Ú!�����+˃��H�S�Zt�HQ�='�I<���)�x��!t�_�����wL��k��~��/6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G'9�и��{4hz�<Ρa�E�Rq���my$�N��o�/���;�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#"0ϸ���f=�NϤ#0��R�u��r��;�~��-�f����Ga�߈.m��B��+�T[nHN��R��bP�63Z�t�5ߧE4��Fr��j�:����|_e=���sg�*��N�{1+�줥G7Q�w�D�o�16�
�b�����ԍk:��+�4������1���9�v_-��\z9ʔsbbj�i0���QgD�4��|���0N��Ӯ��N���E@4"��Sm[o��
����8��"���O^��;M70y���߬�K�"�ޭ;��G�09E�A|���/$�ߺ��]ݸVeXQ��;Әa_�Q��4�Vb6����4��W&��M�φ��<�6�@a� ���N��ȥ�n4s1��7�癆cgQw�c4~Nr_�mS8<�nhDJ��3λe�9�Č��nF���<�W�.�P�	��
�Q�}�}��C˥�!��_�*9 ��b+}y[�k��^�1��dc�@c�����h��-�����Zj���
��I����`(>�������ݚ�Н�;[�T����kb- m޺�����9�q��Ɨs�d�tuѩT��Z|�F�̃��Hd�=ey+�8�Ȼ1��Rޡ�S)W�cМ�}Dq�f��&�(5�;2���+1�;�.��1��!*��*8��!�qgy�`��vN�[���}��4N�J�ף�a�	�+4D@�ݚ�Н�;[�T����kb- m޺P��l_��H!�`�(i3���3rn<F�ڴd0��d����"��
��h�/�f��h��|�����!�`�(i3���3rn<F�ڴdƍ2���l���Ě����E�i�m}6O�D mWN��ܐ�}�-��cR�O�z�U����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ܝ�s2���lI�k4.��7�t�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�TM�a��G��P����U��)���Y;e�iK!���d.���+�^n=\f�5>���௧��T×r���"sS<�0�zG�������&G��������O=�W��E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv����q�D�-c[����dN�<@Iv��nt=:��:5A��p���KL���>Ht�u�UG��Hb� h�ҩ����q�D�-c[����ӲY����&
@!˥�I:��q��k��^�1s�Uo���03�� <I�����&G�����$ZtgQ�9OZ�s:�8���Ӫ�Ġ�9�C�s�4՝� s�#�,��&5d�:�.�N�Ĺ�Z<��A!��-�����d�tuѽ3y��;��"?��FZ� d�!y�b�G2fĉ>99��j���Gp��Ě���aT��3G�IX0F�M�27���^��~"�KT��+Y�6R��M�,!hޖ�A$�P������5d��n4s1�U��B��-��8�2W6��v�����r$ɓǃl[�Ƶ�1tSjv�� �@[�鋽C�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩξK�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�irD3w��'��a��o���H�RtV�^$����}��*�f;��}Dq�f��5ߧE4��;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���r5�I��drB�WD�{����0��e���F�&�?\MP!� u��r��J>zߋ��>ַ�����ƍ2���l���Ě����E�i�m}6O�D mWN��ܐ�}���$�uG�N6-	��6<���oA�LD!�GkǤ661��������C7@�����hH��6�3��N�߿�wW��ZN����6�o8:4�I���c�90��G��6�iI9�o«IX0F�Ms�Uo���ci���{2�'ž1�|�'����u��r�吆v��7�tG��!̒j���b+}y[�k��^�1��dc�@c�����h��-������Ϟ4�>Ht�u�U%��v��;�jmT�#�0M�Ŷ�Eʨ�`N/�a�	�Z����ڎC�?�& @=F�S���iﳣ�N���V�Ո���߿�wW������4Yz����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�m`����Z��b���Q>�<��#b�8��B�5�¹�*��a"N����#�T������oj������ZN����6�o8:4�I���c�90��G��6�iI9�o«IX0F�Ms�Uo����=Djw�9�xjzӝ���I(͂��-������Ϟ4
T�W��%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<Dw\����ō܈��VW �+��}Dq�f�����,����0�|섃Va�irƦo�
�ƳI�^$D���5i�a�vb�(���27:�������&2��OY�J�M����!�`�(i3s�Uo���[;\v�a���?D�8����Ě����E�i�m}6O�D mWN��ܐ�}ĚȜ��Y���܆��줬;}it���U�R'�˴$�#��Q1�dfC0o�4��F�悠A�,��b
�C�&`�@|�v��������U�Rdd@��2�M�,!hޖ�A$�P������5d��n4s1�U��B��-
r�	O)�A�IS���=Djw�9�xjzӝ���I(͂��-����w-)Sz�M�:�.�N�ĽC�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ���U�R^p���P#%��v��;�jmT�#�0M�Ŷ�Eʨ�`N/�a�	�Z���Lm�<o��!\��� fa�н(�P"G�wk���zܳX�P��%�©��-/a8X�o|3bK�����`���UK�"��ӌ�rHN��R��bP�63Z�t�5ߧE4��Fr��jlk�p�+N᢯��0��ĥ�A�)�'� o�F��(�[�o��_�Rv�䩲$��8��I�:Fa�7��׏�������u��0C�r$ɓǃl[�Ƶ�1tSjv�ٮOS���p�]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����-����;�jmT�#*��m�vэ%�K��^/p#��I2�8��[�@��W��*����!�`�(i3,��B�u���Ӹ?]qt���-����!�`�(i3��S�V� h�\��;�,�Ra])n#���r������!���Ĺ�J�E]�?-O딈pᜯ}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��{+�t��Rz�R�k��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�sݸ�/�gxjzӝ���I(͂��-�����d�D��^օ?D^���k��^�1��dc�@c�����h��-����pT/�GS�~�+yp�l�����z����-����;�jmT�#<��4�e�AԢ�a\�2}$#h6��8{4����g�B� �b��!�`�(i3�j<��?����"���w�w:�!�`�(i3u�st�⫴�IV�*F/��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��̓-���.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc63ͼ�a+��X�\�[2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�"�_�Ȫ��q;�4���W�&]�6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&GZ��JP��V��#��6x����E2b�z'hۉ)��d�7�q�e�OB]�4<W��Q��ic)�̩ƍ2���l�;Tti�����|�g�'DV���b�z'hۉ)��d�7�qĝÜ�f��E�h�b��0S^Գ3���ƍ2���l�����g�Z��3��a���!@�f")u��r���\!�U,ܓh�,��R��3��
�M����d��-��!�"ǉ�t������z����-����H������N��������;q5�y�����ݚ�Н��s]��z��(ǝ��� ���c��9��'���t����}�}!�#�b�	����
/���p�j^!�� �!�`�(i3��WDChFb&N"3A�NO��J5�,�Mpf��fĉ>99��A0ok�����F��O�<��}�u嶫IX0F�M,�E�ϣ%� գ>4�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������L�Y&�(G?� 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc,I���HG�G�_O���U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&GK��ft���-:��;��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r���\!�U,ܓh�,��R��3��
�M����d��-��!g��J�s��z�
1���;#o�]�ʄ�v�4�?zm[���*��-����P#+_]ݱ�t�UW���.��)��{.��V޶�Z2�k��^�1��[��o}��MX�w����D����K�f�1tSjv�K��ft���-:��;P�(,�Ȓy:�1^0lfHN��R��bP�63Z�t�5ߧE4��Fr��j#k
z��k��Q�a!7g����]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�x�\o@���T��.��p�캁Y2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���m�(��WDChFbM�,!hޖ�A$�P������5d��n4s1��7�癆cgQw�c4~Nr_�mS8<�n��=����t��{y�mV8��0��1�"��b+}y[�k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vN�[���}��4N�J�ף������&G�B�'��a���{y�mV8��0��1�"�"��K�w(T"c!s��̢k���
�I�8����q �H�%��ZtV1{,�m�ښ�-����P#+_]ݱ�m�
���nGW�:!�EҰ�WDChFb�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b׏������{y�mV8�	՚�^��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������]މ�;�Gۍq��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!@+�ϕ���q��B�`�J�ɉ�z=� ���ɡgJ��E&(p�
�Eu�J�?Ig�(��9��ᩃ	tN�\c�-2���S&ϊ�;ѩ�E��p��u��.t�=EpH��j��A�0: ��q����%	�3)���C*4��]���
@�i��g�?�d���&�V��o5]�:�b��t.�C��6�o8:4ښ�*jl���C>��ӚH�RtV�^����Y�z0=�_���{_8�Y��=�}�Vݨ��}Dq�f��R'cf��>��YfG��-}RY
xǍ�J�r��ps��u1,����Uh1�[��(��;�jmT�#PB��/���߰�$|�Pu��r��;�jmT�#��	�DůI�߷�c/��-����!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H��Ⱥ�Q���'g`$�YD ��� ��?D�8�鉅�%>�rGO�D mWN՝� s�#���k$ �H����ڻ�+���i��ċ�!1tSjv�!�`�(i3
/���p\"�!˥���KS����<;�$��\|����=�'�^�����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��?�JY�)�,�Ջ ��C$�)�vxZ`�b�0P!6j�"Hsކl9�p��e޸XhZ]<�����	��TtU��
g1�MVjg[؎��&���.ԥZs33� �=X����\�5�O�%E#P'}�\$I�}!�#�bM�,!h�z���#A�}?ɝ͇@���8-|�D�7��aM*:�b��t�l��p�xB�my$�N��o�/���;�SENan&�� ���� �KS���*�oF���cԱn�+|�[Xs�g��������:=�)��S�2�]�Q$iP����p��ݚ�Н�X19�-.|}��FL��G��Hb� h�ҩι�+�t2�c�^[v�5�ܾ��mk�9$[{^+#y��MxOܳ����|e"fĉ>99��A0ok�Ra])n#���r�����Jo���j� ��7P��'����u��r��!�`�(i3����Y̀�3#O�2�B���s�����X�X���`��,n��뾦�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�fF�5.]���E�i�m}6߸��S�Ȍ��9�ڮW;��|Bΐߧ �l�}!�#�b�$2j�K_ryQ�j6�S�z�����F�t�ϛ�c�.[K��mZ�'����Z�G�a}C��B�No
/���p�U�.��k��~��/6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r��;�ƽ�/��e޸XhZ����xO<�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H����D3w��'��b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����,:&Ȍ�g�F��6&�U��f�!�`�(i3<���d1x��r-�T�����+v0: ��q�e>%����T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH:�b��tv|	C���0: ��q˕��h `��;b�-�2��;�P�t�5m�ڨ�hծ��Ě���aT��3G�IX0F�M����Y�)en7�4_&��,2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$�/T�!�'��񫯃���{S�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�܅��6���+""�?��n��J�
����[2BĊB�#y�/&*�vW(�����bʚ���"�Ag����<v�Y\`���8-|�D b��tY������`��nF���<�W�.�P�	��
�Q�}�R'cf��!sR*��d�(���B���o��+eQL�0� [�3	�o�{�p�l�~�Q?M8�f2]�Q�&��H'o�a8�J�M����!�`�(i3i}B2>�~ �<j�"�AM?��y�!�`�(i3ʲ��U�4f�
"_��P��]�/F��?D�8��	��x��ݚ�Н� b��tY�0�����V	����/��kOTfĉ>99��A0ok��$f��_Ub��7��G_��Ct�w#��@\E�W��4b��Q+��
���t��{Ck	��+�a޵��	��!�2��\HuE�x�n���R����!k����@�=GGφ��<�6�@a� ��fFMqlg{y����i�q,?5q�D�E���'���A)�'ž1�|�'����u��r���<��a�X�r��ڵ�r)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����D3w��'��b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����,:&Ȍ�g�F��6&�U��f�!�`�(i3;s�e�$X�}���钝���3�#��}Dq�f�m��;���1&��*�("��X2��4�j:��e+�������� h�ҩ��m��
��>W�~����2�I�b	�fƏ���%>�rGO�D mWN��Ě���aT��3G�IX0F�M�~�eW�Ae��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!�0���ɵx�/.ؘ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc6^-Yu��_;��up�6��o�
w�f�:"�G�}��d���!i��f�,�k]�Ǩ����)P<�ܓ�Yw�R���y>��yСs$8��ѡ�X��B���Fkbҝ��q8h�9MHH�7ḩ��H�V���羹���-oF����7Î�I&ۛ��*ަlCi�n�&��;H��I]h���R]�yRy���4𢜋� �^H�^���H> ��݇+�� z�P��	���QC�íN=]b~*��s�φ��<�6�jdƇ�n!+U:R�;�90� �p��w�� ��(���27:�������&YG*�ctB�1����2��wl53�e�'{w#/ B!�`�(i3}Y;�jn�.�g3Zv���� ���Fkbҝ��Q>�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc4�`�(H��L����M�,!hޖ�A$�P������5d��n4s1�U��B��-_S���\��uW������r$ɓǃl[�Ƶ�1tSjv�t�R!ME�'�^��������@|����^a�nu4Bޗ��jw�	���|#HK���4Y{]$�AՁ_�mS8<�n�ݚ�Н���Q7lY��)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b����A�ձ^�Qb�Upq���!���_2��VU(��z�j�Aa�R�