��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω� C�`N��D���ÿ0�^��p�5�
�V���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:��9M��K�:R��,1E�I�?g�f��r�F�5��I^ξ��ݴg��S�ZC�~y��ϼ/U���T���딣0&_���X0���2|	p��rw@	@us�犕/�h����
ۍ���yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-��Yk"1/|sL'���oֲ󄰊־���1N<��;���u��w)�S��X3����~篟|���zn�����f��8�:r&@1�+Q�<�pQ��G�7��kRG��5`xt��R� ��\}Z35�Ջ��D���Ʒ�����ݾu�y+��T����5yi���FnBƕH�N�4�T���±�h�Џ�q�G����\�4�sP	�b\qB��������"^Y怄����v�~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��E_00���/��aG�k�8���҆�|n���:�o�E������G��F��=��J�Й�m����ǥ�P+<�F�z'�_��z�Ӧ�'�b+aQ�wT�	$~j�u?a'���]����Ϭ	N*�b��n.�G�@���y{��O2��@����ا�k�8���҆�|n����{y��J� V�9+�fs �9p�J�Й�m�K�ţoAE�{<��hr�O��C��0��t�z����!�S�?|	���u��u���;�z-�~	2�O������|�OA�
܊��?Y2���3")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ����±�h�s�JFAa��Bzb;ym��+r��JʅqNA��d��1�:�Ω��
�/�r��]���P��`�.�D���J7"�4d�{!o�ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l�����������f���Ӿ���	���q��q�©������5X�/x��-w}�~������:�>:��ʦ,\ަ�It�k\,آ(&l������ nU�IÙ=�H*.�PS���;-;*�7��ʐx�?�Z�>)��`�U+�PAY�b>bb��:
 |ϯ�JHn��z���z�O҈�]V�H7'�R�^Ƒ��,ԯ���gn��Ab�%^�v�yx8�y�5��Dz���Q�^�y�zL͊�q����S��o��հ���*!�ha��_�Ze�t�TWm������L��BqN!Њ��#�ڊ<?@��[	J��;ι��QG�����U�����+�J��U<o^.K�}��HwL�X������VǛHO��E=]A��O�T=�4e=��-?�(�����I<��fҾ��9�Ǿ��q��w�R̶����}͟PP��Z鎬����
C��8q��f�kN�ı&l����Rʐ���zF�r�f�t��6��	���`y����ꢤ�OgZ)[���F�]2�y�Z鎬����
C��8q��f�kN�ı&l������\�*P�I7��-5��6��	���`y���J�۪�'F&�>BH<M�z�]�!����M[��Ǣ�:��6�J�ҋX����>��l%i�-�|�)՜�4��{l�f|�(0̈��N�faՊJ�e:[e��mea�8���B����g��Tݭ�EB�ڴ&�Gd��,M� ?ҡ���y�E�nwE��S��}|��XH�����,>$+W��� j�(����5�?�J�Ń��ɖ�2i�螘c&�'�᫆�zy�g���+
���C�gAO��ً�}�Y�ןw�8���/����Z1`� k�|6�8W�"���1���g�,P�n^P��:w�(�����@^7&ģM�)sWmyY��!둿8(?�3���Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX�����/��&��e��Ӄ�WUk/y@)��u�h踫g(�r� k�|6�8����^�^P��:w���@c
�}�
�?�k {P@2���e��Ӄ�~�k�l_�]��)��� � �����p>��u��>п�p=	�˳͠m�xW��9u$d9��}ϔ���3;�i��R�^Ƒ����"X��[��Q[R�7��z�h��4f��Ԝ�]����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���j�|�{'�8���"�-[�x�X���z��N��ξ������ei4����/����DP֞ �|p�2D:^�Ͱ��Le�2l��4��a��se�ξ������ei�^���?�������bpP�ԙ����X�/R��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX��}�
�?��+?B�OAW���D��g����H���	N^�U{xN��i>r�<Uee�,�Aٺ�Hr7O�j��I��'�����3ml��nL�,�7�ܥ��2�
������ǛHO��Er�H�8���#:)NV�A���rX� �G ���9��c��Yr�o
�V�6IWJE��=E��:���U_�+X�V�0F�Z��cfo�*�Y�E1� ��C�8�J�Q������2aȟ�h~��b!��uፀ;��tJ������XIb�(RzHS�&�h��=���{lGD�V�B��иܖ��A�.u�rc⽣�Q��'2!2�X 37�˱�5_=���$�4�\_�=@�G���r�ϸ��#|ShI�ˋ���Mei|��sD�hV�\w�4�	H/�"�����ʛ�M>#�!�`�(i3Y%T��BP��&��J�UG�s���#�n�%�y!����-!�`�(i3�a�\����8x<�A!s���Z����Xc����L�{Y%T��BP��&��J��\��;�,S:H��+܆} �S�
â!�`�(i37�ܥ��2�A�Jr���CVF��g�M��p|�\m���X����)�ak�m6���D	��U�l>o��|���bǬ�=����������622��fH��>d]=]A��O�T=�4e=��-Y�VN�=�ԃt����}ꇐ�622��fH��>d]���+�J��U<o^.K�}/��<Ӭ�/�"����J^L���I�PD�naзq8�Ј)w�<�_N`E�cvR+��}Dq�f�(����O��9�JzM�E����F���8�TP��@E�`�8���&��#�@�o0�&�v�x"�,�>E��ʆ�In��tT?�7G|`Y��j3��� Q�N��*lOO_NK8��40=�4e=��-V�׍A���}Dq�f���<E�f��V�mK�b���G(������8�TPO������=��w�[�4�Mei|���)C1Ew\w�4�	H/�"����0�:C&e�!�`�(i3!�`�(i3�a�\����8x<�A!/�"����kU0F�o!�`�(i3!�`�(i3�a�\����8x<�A!s���Z����X�B�r��!�`�(i3�a�\����H�:"�\�(�6k�4d�����͈��}���i!�`�(i37�ܥ��2���kܪ���*�LNm�Zt%��m&<2O!j����x��B5�!�`�(i3x�]�V���M�K�=g�H{g�q��������b�Xϋ?@,�Xʚ@h"�,�>E��4];ˍH��!�,���;���2[����|��1���Wʁ���p�B�E�!�`�(i3���+�J��U<o^.K�}/��<Ӭ�(�6k�4d������z!�
�W@!�`�(i37�ܥ��2�`e7��9��×�>�濖��#�(y��K����!�`�(i3�E����F���8�TPm=_g}b��t�����ܗ�J���� ��A?Љ'�-o��`%��)w�<�_N��M��+?���C&��>k0��w�*�fBg�!�`�(i3���+�J��U<o^.K�}�d	c�b��8���&�Q�$_���]��3a��!�`�(i3=]A��O�T=�4e=��-Y�VN�=��`
 ֢����e���W��]��3a��!�`�(i3x�]�V���t�����[F�a�+�6�5�p����Rܖ���B�r��зq8�Ј)w�<�_N`E�cvR+��}Dq�f�(����O��]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=~�Y���(���8���VZ��W�d�"�,�>E��ʆ�In��tT?�7G|`Y��j3��� Q�N��*lOO_N-�4��j4];ˍH��E�(��<���A�� ,�ttT�r�pΚ�w] n2ϒ��[����r-����8�TPO������=��Z��( ���~*񇦳��Hw�6ٿ����зq8�Ј)w�<�_N�b���VVA�ڦ�c4���ɺ�y��k��)0��=M��LO�|43��52נ޼��X�B��+ H!�`�(i3�E����F���8�TP�}O�6`-�b��Χ�����BQ�.�`��SxEWI�I+�!�`�(i3!�`�(i3"�,�>E��ʆ�In��t�hFyu�.��J��ߟ{�����8n%d��z��BB���#��`'��e�x�]�V���n:�t�c{DJX</��}Dq�f��D��[�
�:�I���G!�`�(i3!�`�(i3=]A��O�T=�4e=��-�ĕ|G���t����}�[V�ct�!�`�(i3!�`�(i3!�`�(i37�ܥ��2�A�Jr�۞��Ѵ���t����}�-O�9�nd_p.���R`!�`�(i3!�`�(i37�ܥ��2�A�Jr�۞��Ѵ���V�52SG���C!�ªj��졼�!�`�(i3!�`�(i3�a�\����H�:"�\��|#HK�����\��w��;�����e��H!�`�(i3���D	��U�l>o��|��@	J�!���}Dq�f�!��I\+��M�a5��|���瀆!�`�(i3=]A��O�T=�4e=��-v����]c�VA�ڦ�c4#B��F�7�ܥ��2���C�0��(����r���� �G�|o#/GD@�F��q+�#�!�	U�E~�˲�<�!�d�<6E[�:x��7JS�����,MLG�j�.(Wx*<�6�Q=�;~����%ho����G���r`
 ֢��FE����墝{l�f|�t�K��0�!�`�(i3!�`�(i3!�`�(i3�;C@����3a�LD�P��Μt��/N�M�O�IQ���}/�"����Ʈ芪�x+�o��C!T*p�VU��J!�`�(i3!�`�(i3!�`�(i3"�,�>E���� &N��nF�d����M^�{�W�Q�
_�J�g�J�LQ��w�mK�#]2� r��w��S�)37J*u���{��}!�`�(i3!�`�(i3!�`�(i3�b��1�K�+��o�.@��A�OH��*Z�h�TD��L���2��}��g��9|P��{l�f|��rs�i���YN���G����exa(􆿳�xE�zH^�7�{_8�Y���˂lq�㜯}Dq�f�F�d�����r<K���J�LQ��wEOJ�uxm� r��w��S�)37J*uc�A�L'�t�O#��XvU(�8���/��}�Ш���my$�N��;� ��b�� л�w-H�.E�^��\=��
i�c�r׽v1a{J�:�r�7��'���Xw�j�7���N�v�1�����7����`y���ȓM�Me����Μt�'�al��p��B�NoSƏw0���8��Q<��z��}�0z�cUL��լ[po�uYG*٦� 7�v�ԯ����fbK7͍��ճ��)�ȓM�Me���섫�So#�'�al��pz��+��ݘ<�6�Q=��f������L�}*2#ԷN�ڿy?"S���0S&",f�e�0�؍�3Ϟ��M�+,[�� л� Ƞ?�T8�� л��d�Q���S�"���=�R���=�u@Ý��},��X:���v�,,�kQ�Ǐ˨�g����K���=
��P��bE˧�<vr/��S�s~�k<����-Ի�弳$��P�!Ўx���-�z%8;����v{:��h���1���N��X�'�f�E�k�8�"�$�����o�u�/z�u #��Mgs�4�H�O��	�� ��Fw"��Aњ��f��>�%Mg�� л�G/1avQ�e�b�����,��Z?m��r�գ���VRj8�@ʚ��X��9�����Ïb�}������c�.D�"]�ϓM���o��C!T*p�VU��Jp��T�����hy�%���[��S�)37J*u�,�JL���*��c�d}];�SS�qL�\�Q���}�+�^@��#	Ͼ7�Z#^L�)�4)	���E}];�SS_�⥳�"_!�`�(i3!�`�(i3�� л��У��a�p�탯;\߰ �Ye�]r��8���F{�grT�i`YS���UP��v��!�`�(i3!�`�(i3<�6�Q=�U�"���M]�B��5.��$�]��tK�"8�f��>�%MgY��j3���d=���ǄҋX����L$�����/���NM����s�٩��8bq�Be��]�!��5��E0�ƺ'���g�{ ,Cѣj�k�-U�P�d���0\��1���FM��`��\n$̱~"��>d�c#�'����1���<��$��tf�E�k�8�"�$�����o�u�/L=x��gO�+�-���qJ�?�̿��{Z�|bQ��� Ǐ˨�g����K���=
��P��bE˧�<vr0�����i�é�I���z�S�*��iMOPԙza��5N�ʡV�l��� л�/�ދ}Ղ�� л��d�Q���S�"���=��
��L����1��in���� zԻ�弳$_N� ���ui�X\�̈́nlH�I<�6�Q=�w�3����f
�@"��g�����R��H�O��	�d[��K�pHj�4�\��ލRC�|�"u�ۼMQNv�2�^��)('���Xw�����C���������C���/S�)37J*u�,�JL���毘3)�:�6�5�p��nz�����:�r�7��'���Xw�����C�������ڥ9��[ʫZN��ҋX����L$�����/�����zQ�.�`��Sy2�H	�?��ҋX������S8��=�I�`A��8���1�pp���aa(􆿳�tP"7��%e��0�U�S{����<�6�Q=$�D5�bY[�q��7-]P2<WV��
i�c�r�(����O�����b3�'���Xw�j�7��$�~����$�⹌y�S�UE^����Cҷ��e�ˇ�h����2�[Q	��
�Q�}#�ҒIs{S�>��{A��"�����f��z�� л��Ujc(h�t�%ho����G���r(�:�f,��iQ��e�Z鎬�������(����} "m��^�V]��}Г����ѓ�1���`���A�O
i�c�r׶|�ل�\I��w��,c�A�L'�t�O#��XvU(�8���/�7��I+�:����fSM0.��4;�. ��F����U�e	�K~9M4�6@|�y������-&�6��_���9�����d�J��:�����"���혅vº�w�⽒���M��ҹf�f3';��|B���r����~?ш|��U��)���Y;e�iK!���d.[�����:Fa�7���^�#�n��Hc������l��A(�c���_G��Hb� h�ҩ�?V��j�c���o���T�{_8�Y��=�}�Vݨ��}Dq�f��k��^�1��dc�@c�����h��-����!�`�(i3e<�Ia��la��o���H�RtV�^�2��}��1�O�ᬧ��q�}��Ps���'!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�ȌW�7Q�ǭ��w&�.�V��	��y��k'�Q�1\�7� ĂV��	��y�v�g ��#4T��d��Q١Ӿ�$eCD5�*
�5��Dz�ͽ?ڄ��5�O�%E#P�� ߌ��9f2Pih{���N��w
6j�"Hs����q���ط|����B�x��?�_V�VG�88�;矷��N�����?�d���&�AYA@�� ����^���uS �����I\��!��6j�"Hs�x[����k�UH|�b"�uQ��z/�B{�o
�s��$�Z;��|B����ɠ�o�'�/��T�lw�_:3w�⽒���M��ҹf�f3';��|B�V���p�f�N�<�e�S��?�F�^C��}�t�iZ]XF�hx��G��!�`�(i3`�s$����j���9����������"��O�9��~�90)�ʆ�In��t5�	�3)i�?�P����f����6��ͯ�����3m^�ۘ�}�ɶ��!�`�(i36���GԸ�����k S���zǣ©����0�C�D^J����'�kf�<�I�֐`�A^�!�`�(i3�+�H>�?ۭ�����bJ�]�R�r�j�b#!�`�(i3�+�H>�?ۍ?i���7�J�]�RU�`���!�`�(i3Y�b>bb�D���;r����l����F[`3*�!���6%�a`�3J�V�h7�mEoxT2`$x�������� Ԝ93����!�`�(i3�q��&�X�!�`�(i3�)ύ^��R�^Ƒ��f�?ǉ�=��x��&^]?x�v��X;p`�;-;*�7��8���168ORN�]�5'�ݚ�Н��dv��oTN֢&@��&<�6�Q=����@4�0 L?�p���@ZZt%��m&<g+b󆤐=�0��"��S8���#�j[�j}��YF�����Tg9��!�`�(i3��#6q�Tl�������l6�Y��j3���������g�Hn7�(�!�`�(i3��O�q�̍YY~����V�my$�N�����Vx!�`�(i3HCr�1�s������J]z=2�4��*L: �i!�`�(i3�֠��������,�ǰ�m'�2�ɹe�fwy�6j�"Hsi��׷l�mp��'�V��rU�w�⽒��8�>r&�,�Aٺ�H�f>x�:	�W+��W�A�~����Ձ�=�n�V���<XR�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P���Mڷ���o��[u/̉�#��_�R̶����?Y[#g��}�	76�&�;��|B4<d��
~�{�Bͳ��;��|B31F��~Gf��x��9�Mgw�� 
~�F�,���XF:��GZ>.�0����ڀS��d���!i��x��=;Y�ۺ�Ub�!�V��u�ct�:��REs�N
�u�}�T�\ ��;��|B���r����+�uB;y�XNAA���v{��lw	+z��D�H�}�	76�&�;��|B�T'[/Ʊ�&UX�{6j�"Hs|��^�p!��y�;�{(㷾���G���Ld�-P�Z:�E����FQ��ݢ^�A԰�N�5Nleo�c�0gѷ�/_>�LD� �B�S|�P�DM몴PBoT�R�f�~��(�
t��Y�{'%s�Ǹ2����E�vwx�k�g��U-�enzJX��o?��K�U��]�!��ߞ��-���o4Î87V<��z��}��@5���<���q?����OEǄ���]�!��	Ǹ�y85��3}�@�7��?E/6Ұ��8_�����-U ����q?��0ǽi�*��]�!��	Ǹ�y85��3}�@�7��?E/6 K	����n����-U �j�i�K�A��o��C!T*�q���U��E��v��])���/�Z鎬�������(����c�<Q[j��"X��[h<��BSbD�L�x8��E�6ɀS������FQ��ݢGJ��AK �_"p��W�W��<��W{0`�A1�2Y�a��bft��N���m��;���g��I�|�	̍�������������p���Ї�J}��M^���B1��?t7u�`'s^��>\{Ф�E�+��c�4];ˍH���@E�`+�8�lc�@hG�������p���Ї�J}���������O�G��o��s4k�r�j�b#������So-�>�6C�(�HB���ګ7J��n�1��ņ�}h$�ɹ��I���x:����aR��W��90E����4������y�;���g���W��90E����4���"5���q�؅��FJ��/��<Ӭ��W��90�EF�]�`�|��K�z�ix	��GD@�F��q��M��+?��>�F ��>��d��vVx�]�V��v��K.Ū��lEs�/@0e��!�8ߗ:w��y�~��ۢ����ˢI"5;�:�=�pY�~ȸDz�b9����$�n�������=YU�p��.��6ǿv�ɢ������=���a��z>�n�S���=YU�p��.��6ǿ}�(C#ƀ��=���a}����|��t��o�5!.��@h�^x�]�V���\B������d�[�[�_���勤U�@k����c�Zw|�pMGD@�F��qX�ʟ��{ŌX��V�t(]�XnS��z��`��
e�$j�U� ���_V�׍A��]tn1\���w��-��3O�v�ɢ������=���a�`��	4Ij]�������Kߞ������|�7����s�ݺᣄ�I^Ɍئ+�����R�:�%��X�B�l�2�vD���?a@!~�X����Ѵ���4�H��ZX4�x#$* Q��Esȸ�"rR�����P5�D������o!�� U��!�`�(i3���+�J��U<o^.K�}��2����p��I�=�>ll��4?��X9���		���@!�`�(i3!�`�(i3JHn��z��r9�3���Fz�Y�b>bb�D���;r�!�`�(i3!�`�(i3�Q�^�y�zL͊�q�����7�f�ޥ0D���>M�J<0L}�U��!�`�(i3!�`�(i3l0��F��j �i7�sp>�(��&��Rm��e��Q�Ȗ~B��?�d��!�`�(i3"�,�>E��4];ˍH��\B������d�[�[�_!�`�(i3�*���<�Hr�»�>��-U�f��Q��z�n��!�=�4e=��-	i�/B�6��&�eP/�1�w�!�`�(i3���4����4Ieŉh!�`�(i3!�`�(i3%Ah�%4
>��XP���?W��q:�5¥������c�4��s�_oWKP!�`�(i3!�`�(i3JHn��z�w٩L7��!�`�(i3��E.t�