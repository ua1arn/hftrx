��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#��qK&�+K�����Ӑoe[��p�)
ARa��]�5�6�0��c�L��k77Sp����"ݤ�O�B���dW��mx=��������@^�!��s{_꥜��
��k,"��s��)"� 8b@�5�@4:���aD�����9���1����-cD��a��?�MB(< ��3�x �9�T;A���=[��4�16 ����ʔS���C�p�\ �ý��$ƌ֯���.�抳�����y[�39Ye:�J�o�1R���W�/!����	8�! %Zy��iMA�:���m�a�j~"2O0'Uڮ����_�c-��A�3��=�.c�`3�vLC�>�)'��I�����������ɖ�:9b�]��GU �&��2"�t�$�����
_��{T�����G0�8ya%q�R���a�ȤȠ�՟)��+=��{�d�޻ݙ��o�Q%��u=M�q�yk���M��.-]'�?1�z�T�O�τ�r#P���^-�P�f����+�+ҊMsK�ָ��	/�]J�2>ը��;��m�ˋ�ɬA��)�z/J��rH݌x!_w�a��Q�{-������o�,�7n��g\<��/1��]��N)�gY&�@���/�&��z��`o%:���ư����5Oy_���gr2\�D�Pd(��k| �;��f��Qkv����B�Mɾ)����M9�_��$�"�
�I��0?��
+�-5�l� �`�k�ؠ%�z�$�p=�K���� ���;���K�
x���	zy"�O\��@��N�������� c��ǲ����_�ؑ㧝U@�x��:=Vީ������<sA$�v�D��>�����Y�R�[��s�x}��s�7����������X��yc��SG_X�oi�ʏ��~B����R��x��ߋb`�Eın�l �_eS�l6�_1'h2N��[�X���uu�Ǯwx���%�2�/������1N�jAy����ߟE��^7Ldؘٙ�^�_��Xѝ����D�G�;�Ś�YJ?��vX�"�`�/���:�+�Mhѣ�	�J#Њ~�E�cg@���X9�^t,���H�l�'���+�=�ג��S@�k�N�� �m�2��-5?�r�o�ӌS7Ro�Q�S��+(���]`$R:Dza,@�N�?'�1w6SkG�5qv{��Ɗx��8�9~X��E� ���TŎ�ɯ�[@F#x~����±�[����m0�ҁ���)Cmr���`0��oS�Ɵ�3�~#	����Qm�ը����c�)��*h碫���h�$������$a�W��+�m�j��Ӓd�c��m@���k�P�3$.�ǽ�M�Z�ShF�qK}��-�G�{�a���z-��gubܪ��D�}�ny��v	�MLR�Pa'�K����d,zy�I��v]�܂9��Pׁrk�j%�V��̭�N!W`i8 ��XrZKTb���Q��=���~O���/G�F�ՠ�ˬ�ZIl��|Za�D���+ֆ�$E�o�����w�=nZȖ�/ށ�e0�@l86'����L�<>�p�� ظ}J�Ȣ�D�d�c��^�S�9��I^�ڤ���̗0r��з�L�Ȣ��$g�3[�X��Q8,��d�F�"fRAnT�$T�%ѳ�C;^�8:�5T�ԥL.�T<�{�3��</�-�״�.:���3y���׭�����j�YO#����ӯL�aD��ﵵBxg����ř^���H�b�vݤ"?@���7�W)K`'��������}s2�@�!�����[]$�zJ��L߯�O�G�w���'�@H]���g(������@R��d�iLFz�u��YPDv~ǜ�}zι��-�B	]�`�<c'P�Ǳ^\cuO��+�6�+`��c���Ls�O܍��Y�M Ө`�+��T��+��*��i���"`&<�	���o�����~˦��C���*|�ȕW_�'�3�)���������!�/0�#�,�Mp�~uݟ���<��B���d���@4��o����G�Í�P"�A�o[ef�I����4��j�Z�`H�������ň#:�2d���r��(+}U������S�����)�G@��k|�����a�LŁe���8 $t2	3�cK��wa!��#w�H 8Nߍ��y,��u�L/���oN�(�G�w3�7�z9 p���o�35D�[�F�(�倏�5�^�OԓM3=	�0pӍ�@�Y���]���ѷŭnC��l}�G���P&���5�{�XtdP,s)�N�_�d:r�>A�FMWn8���F��ӈeE��&�.��ELz�p%p���n)K$aQ��ج_�Z�Q@�ͪ�y��Xb�џb���˵r�>��.%��yt�Bd����'.�2`�?�V��	ls�=���W=�xR+�t�ݔp����\W1��M��T�0�T/��.�2�m����r��n��ݲ����zl"��	�e�wT#B4l���w�@���?�9(��=6�e{�z�V(���?����͆Q���"��KMVXT�d �0|^�@s�������
*Dz��RذP1�����f�f*�W�d��1O��:\𦉘� ��W �����I9j_�vV�{��+�4S��	A�Ps��$j���`h��F}���2��m`}�-`�F���@���~X���j�8$)�T���Q<)u��xw����˔�̌��޸%=�󶔰��޽�_}.�)_)%��c�q/��y4���)ǜ�<=t�Sf�����3���1��Kb�q�K��[#K(t�|��M�����8�d;X ��m��!D�qJw�xT��k�