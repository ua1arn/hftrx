��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0T)~�������GG�Y��>�RK1��i4����T�d�W;�IL1_��F���֠�,��&5�{�
�<��F�FI�6������M�wA��j����nD�Jy�f���1��q[u�'G�׫� 7�V|TT���B�K��xi�]0��Jl��,ٖ���wL�AZ� ����N��,���m�S�&jJڽ���]e�����.�a) �Y��Ѡ�� *�G�$��vr�[����W8.�t�}֘A�ۋV��J�U�s�1[��Ω���eN;)Ǽ8��s��d��d�5uC%�W�)h�b����;�!k/>{d�'�o�H�{=֯+5Y!L q�Z�&��B^_�Bk���b%�#�����-�uV�"��ą����mѽ��6b�X9da�S������4���oh��ǟ���綞]��t�ݧpUv�S�^t[�0ꀬp�~�Q,������Es0�0!���Tu%T ����L�d���Y�f���k���L��B*�}t6b�3�,/嵛�; ��ܕ�J�O�~���˕&_����F0�ұm��9�����8m��	�:����&rh|���E��j��+�I��Px�,�>PU�ǜ�@cM)��Y5���-��6��*O:���Q�W���#:�aδ8��$0�@����Ƿ6����	`k��&�g���@Dr���'��\l���&�<A��
Ğ���O~����XJ�kX��Z��Ļ����o7'�V�r�9\��F^As�u�~_`���X��Ǝ���q)7d5�,R"�ҍ���cZ�eZN�xM�3s0�&&Q�����#����5�W�����p��6��\��g�X�{����l$�	X���4� ĥ�˙�5���!�%K�Ha��T�J��ay�,T��wV~��`R����32:?���Ƙ[J�}q��
���V��*%Ĳ!�Sm�����3 b�IYT���D�;���:֭��c͛��ijS�5_�c\�=q]l&4	�/�o͡SR���3�;�T{��5W��gnyt�G�,w'<���&
��9?a�Y���x�޴�v�=�i�;��+��6�4��)˟���^p(@U��H},.�O���ҳU����e$�{y�@cz`�W�*
^7�'�S�F��Q�"�~E��m���y�խ�uL��p�`�G��`j~
bT����Z�V����������u6�C����3n �ͧ�2F�M�V����3�؟K��w���e��(����$��p���;�Ζk�4Bw�h�}#Z�f����kR���V�[���l2C�q�(�l�`�ݞu�~�k��k�ц�/��P��Z�EdԹn� ��5��8o�<A��%��7G�\�IW�����@Vi��:q�9������:�m��Rk骡�'�r�T��Pq���1��ǹ1�����c���N�(�gAD���Ap�|��N�F6uh���C��x�-g�}K�@AW�,��`���F�������#̴(kl��ݝ�� ��"u ~�Xe�󴘧��$������p?���:��Lj5��/h��o�R���-5�.�qP�p#�&��ǻ.9���6�jN��DteV�a� 82������xsU��iGܔ�	�ע�R~�4%9�wR��&�T���Y��1q���0tӮ�.�D�(^A}Գx��!�,��rJ_��ܤ]_�����2?���&A����x:���W �}�'ʿ���Y;��9:�"���;���P�zG�ڏ"�v���A��al�'��!`���
������	w�)�b�^+�D���A-3p^x�w�\_��d/cL'Է���&���l c���G��^be�W5��|�AS��,�R���Y62C�tw�>�{f�K	�i];��H�{�MG�Yx���r�Q�ܘ����cjǃ�[��$q�b�e�pA��Y�1I�s/�/�m�����w���y��vɺFH��(Hn�gR���0�߇^�頻,�]���P~��9��#r$���(Z���8��`*�|H�Ճ>Ĩ�b���hs^]�&2��w+��HP�N���[����{c�-�pB�]%ϲ�8)AI,��''u0!/l�KT�!;������a�
ý�;��VQ�h{R�I�L0槤�		���M)�Β,Iۙ��8��4��G�봂9iI=��q�Y�ќE#-�P�8b�J>����W�N�F�0�0X�h�[.�"q���9����_2�b��SW�Ƥ�̦�sB_Aj��ź�R�E�b�,y ��R`��`	*&V���X�V��?{�%�b�g~<l�(�Ol]뵹=��l�B�W6.�޳� �J�ԙc��q�f�=�1����U�ݭ�H�� ��<r�:���@��z��] y��:累	׾���g�3�����7��u���(�1�����e���	#I�Q,	���=�)�:h]#qT��q���{cb&�
WW��<�ˣ�;^��]��=~j�ʯ�s�79��� ��IEj���<4���ϣ!,U��+�| f*�jy����%�y�6�,U�9���tO�LҘ ��$���6z%S�H�s�AG��HIGJ��/����N$�9�Y��Ap*���C_�OmT婫�b�����q6vD�rp�����i�jO(�o�3�<���5�W�"��S�J�f�w1Wv�x�����(���-�J��8�e�a83����zW��u},	�����<y�@�5d�N�|T!l���G~��TUYL���O�rWB�_�H&̒ B�����I�/�U�Չw�T<g�	:�4�:l�SƁ�T�8�"(��$�[���{�E\���w���DB���18�=�Sf6�V�ͬټ�Ie<N��ݥ��p8�g9�L��F��Gs��y����o�Y�д&�O91"FiLa��<ֺ���?a�8|�Y;{�c(�G�nl�skŵ�ϡ�h��~JGt�yfX����ft�T��fQS��!�`,�}'�eڛJ�c�1P�N9cJ�]yo �q�`�EK���6a#8b�W�Y�Ch�odQ�=����I���G*��s�Hh���N(A7�h�?���MJ���k�P��r��F��7�Ϟ�V�T�],_������^���G\��v��Q���Mp��N��u��eQЊ��jŠ;7��ҥa�3��'Oۖ�<W���ֆ7�@�?bH���UU���o��6,�Tm����c��+�b�_L�zF��2��=�8�zH��N~��kP��!�0`�v�"@��O�$u�%P�ػ-�Aʁ�ջ��0�y~Ijo�:]�L����,��F��L5����r��_�|+� �To�����g��/���mh��m������H�M�.��nx��}0���X�r�I��:Dbp�|Z0�g������A��a՜�	�8��M���p�W���&KGVX���a6d������`������i��NJxC }��G�$4�K"e�&�Yv3���m��\�B��rA6�?���	pu�p���
�dN8�a�i��K�#1��{��muo?=�����<L4ą��qr;��B�v��R�2T|����5�8rG�%7mj��{-����� ��RmP�ެZ���O���3�/ż?ƚ���f��}��P2�i�T��)�\�x����J+�u�0OJ&��࡞>����f��rf����g��,Cwٹ��_+���i��KM��4���7�����6M�S�MV�^-Zh#�3P�=OKqd�TBj����QS�#���:��ŲCe�@8������vԠZ��d�ӡ��V�֤���ZJԢb_�������r��G���o1����H"Q̲6�!�]�w]r}}��Ƥ��y-��f����}.�&�߉�Ȃ�[5�&���nOT0�,n��p���^w����,ʊ[H
z��*���-B��~�Sa1����a����.h���� t�.,�F?����nB��Yu�����t�h#�+����9otJȺ���t�(�3~"��~Yc,3!I�:����)��P�|HP�y�9,y�Bv�<����ّ�������v��ۂ���q��=:c�6�а3�{[�"<�����P ��ʵnY'�1�)��q}o�uw*�n��k��r&�p������˕D͉� |@,_,*��-��p3�������,!��Vn��\��#8IT�X���������[�i@�G�R�̙h��ZsId�����3	�u�J�z��/=Ԃ�Y���P}�M�&V�U��Ę�p~�#8uշ�V�/��ئ�7��{�k�7k �Ϛ�����	`�<��d�G��"XҕAܠ��-�!����OU��>t�S�fe!I%�2e����Aq9��#x2gZY���Ss�hn�;��_	��0�@}����S�  ��y7�EMb�E~�px�CX�w-
�^�m"�ޢ#����Ia0͆}2�FUHI���4D�j�%��'HB��'i TA�K_��g�	s�8,~U]:��d�c&�}R�Ӌ64F.�,�`�?�̲�ɜ�c��sgf��N*��)�&��.[�B\���w����px'e���^&6==B5t��ao��!����ƿ�S#I�&jf�:t�e��:<^`��
��C��f���㲕;0����i�I�i���a��h���� 6c^��ǐ,f����N�)O��6���
Lܚ�D%�ڬN7ۮ M��)K�/�X�N�lo�������kfPB���]���8�Ī!<�Q+H7����li*����"AR�������"�z;��͗Á�U�V���ǃ{^V~���j��vο,vw�?[$�������|w�B��ūI�kB�{(�.�JWu���@ڗ�_���o2Ͽ֎��p�E����IFx[O�=�����/ϔ�7a��ddM�ȟ��+[Īg��7��}V�����5]���3��593�5H�(���:p8�y@��'��"?�}�4^_1��BZ�E�����;���r��$&<�{�����>��\�m �,3��r���T�f�y?��ФS����~1��n˺)�2�#9��ױh�͸ns�~&C��%� b9d7�/�� \ h�st�57�9
c&*�#�D�E@�z���ɐ�I�ч�Ð��~����0�7�F"TZXe.�*���E��?)Z�ӈ��抻Z')V"��iX*{�9M$�fcWÄ�jG���Y{�(��D�s ��9}�)fx9��j܏L�U(�C<\b$]��,�c�~v��	 �?.@H�v
���ϐ���N�}�����@����)��iXq����.��A>���9�!&F�:�NE�r���%cO�0���d梋�mj|�z�����١5& ��;��ku��S_ĹX�MQڸ�zV�N�f���AŢ@��ݸӏZ�7~IL���-b�zWB�쑴�?��ْ�F��s�[��տ:�8eR���s�X�J��e���'��`�m�W����N�~�ᮣ�Ԉ5fH�T��c<��G%��6Ib�'v�Ky^d%J:z,u+��z�C�tn1�� �V�)��2����D\<a�
u������o�J�A}��PU�V��@�|�_Ǝ��uc�@M{QZ�����􏎞B�B8����䁏��t�Iiv�)g�ꄊ#���� k<wج҂v����ǚt9�Ň���{�c��L{B($�?+[/�Y��	�c�5�lVOt/�B�9���Xo5�GC�*��I�ݒ�	�H"8^�]����W
A;}ں{�(�y5��̳hP	�z��m/�g�,nwi��_J�H���^��v(c��-��0��x��Eq;�D��Ճ���k�<�s����t���?����N�)� ��K�&d�İ~T��67}��ʝ�v����r(�B�I҆��x���� ��'		""�}NS��rh�`Bz�E�%w��E���vϩ������s�'rݓ�i�6_�_Gx�r������%����d�{�P������bY�r��~��� �<�ao��>@��d��!:<��BP�>;�6�/k��;���ŷn�隢�_1�3���%����K8@˥��'� (X����'��L��
2*������9��4i�G�9��~��z�k�R˒j�_%�f�օض������~�G�
������y��rJ9X�-�V��O~,����