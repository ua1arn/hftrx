��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9|[�,HJ
Κ�P/�u�x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`��;�É_g�?�H�.J"����U���T���딣0&_���X0���2|	p��rw@	@us�犕/�h����
ۍ���yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-���m���.GJ����1o���Nx� ���������	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"��-h|,���(����>S��ә�����/�4�}n'���a*�x���� ����ޙB!7����ˉ�1�:�Ω�>���h���|&���ukh��s��v?�%�ea�;y� ����t��A�sxW�O�k�c��`��Z�>)��`�U+�PA����Kp&����-N�ʆ�In��t��Q�]���h�S{�5��lW0�±�sR�{F3�_� ��"����5'C��[����Q�n���{�)w�<�_N���i��I<��fҾ��9�ǈ�5�G
m��u��N��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�D�+���8�<��z��}�0z�cUL�n����4���á�~O�"j���b7���Øfq�\E��0�ŭ�����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��Pc�Xe��TD���rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0���-n�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�eן�-�Q�Z/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�ЂDa��(O�J,���Z鎬����F�71�B��O1��m<S�)37J*u�񁫴}2��:��ӰӒ1�:�Ω�>���h���|&���ukh��8���e2��'�����N<���d�k��Yu>�G Oag�qod�֓��+��T����oGo�Z�K����ހ d���c�u:�^Y;g��4��s;�s��&<�w�п?G��q8h�G[�� 4&Ƒ:2�c<�^<�H�U�YQN`V��	��y��2����8��`+S6E���7-K����}�)��E�d�-���geW���w>��Y��$1&ODQ3�z�sis@�����]���ϸ��#|S������3[�u8�J�a3mPy��>/' k!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�����hWK{m35%7� ��yDg!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����hWK{m35%,�!�H<�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��Q�V!�(�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��%}w�dN�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�t� ��O���}���i!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�$�V��bst�N���!�`�(i3!�`�(i3�X;p`���z�����2� ��=�<���� z!�`�(i3!�`�(i3!�`�(i3�sg]�_�}F�r�f�t��5Z�����N���96!�`�(i3!�`�(i3!�`�(i3���I�=|�0��E|�,���6%�az\�m���Iϕ������z_۬=�!�`�(i3�&8�,�g����=�'�j���#�|M�d�>b�eIG��Q�q>x�-#F\eڲ!�`�(i3!�`�(i3��g��E��� ������$Y� 2��4�b��{�P}�!�`�(i3!�`�(i3�b[�u2�G�=����ڄ���������622���k˗S�d�!�`�(i3!�`�(i3@�C,��ǣ©��S:H��+܆} �S�
â!�`�(i3!�`�(i3-���d	c�b�ǣ©��S:H��+܆��K����!�`�(i3!�`�(i3-���d	c�b�ǣ©���_`Ogkl@`��m'��r�Nt[NzigzA=v)-��,ufOX�mCf�?ǉ�=�$Nx���t��y(�����������(����������)��-�L�߯d�8a,�X����>[H��_0Vձ!�`�(i3!�`�(i3�&8�,�I���Ut�es��O!�`�(i3�N�v�1��B�r��!�`�(i3!�`�(i3�$wq�����0��E|�,���6%�a����>[HÛON�?��!�`�(i3!�`�(i3�&8�,��w�Iſ�Κes��O!�`�(i3k�-i�9~�!�`�(i3!�`�(i3!�`�(i3�u~xgA���������6%�a����>[Hs�?����H�Ud���7!�`�(i3�&8�,�|�1�0j�~�Y���(���8���VZ��W�d�!�`�(i3!�`�(i3��5�q	�`
 ֢����e���W�\�h��&2��>/' k!�`�(i3P*N�2���9�����޲�e S]#�e����kn4@Q�/�!�`�(i3n&����_�a�/!O�f�?ǉ�=��9K��r|%oO���m�
��,!\4L$ֵ���A��)}�����*��hy�t�]�|����*[UxG!�`�(i3N>�X�5G���oy���ݚ�Н��@����MTl�������l6��6�5�p��`�T1)��/Z鎬�������(����z?|��f�?ǉ�=J�a3mPy�D`}Q'���Xw�j�7���z��0��ݚ�Н���O�q�̍YY~����V�my$�N�m��y���wӨj]h��0kI��h��d�)bU/�'5���ĭ�*�����X;p`�Z����c!�`�(i3�%]�N����%ў׫�t�$��o؍��R��w�R���y_Nr`e���4)���>݈��K+:��0	��