��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�
TB�(+�
mQCJX���6��2���;#��9��p�����%7t�p y�ʌ�����h���./�g�q|�&�y��S��Π,�A{�-�p�3������o�^��ޛ�������(]���M ���l��Q%Soά������iw:�Ǝ�i�O�׭����D�ԫ��*~`C.z�a=�=?-L�c��Z�	>Ԭp�
��B�2�T���T��}8���6��T_�ht�9�r�+Uz �ÿ$$��v�������(]����!�|��P�B(��7�\)����4���C�K)����=��C&��f��kՈm;�C�XTg��	���Qu&$��v���J>7��9�J�GL�q-���CpLL�{���]v�o-S�L�8d^���5�WPU�^oj	I��ڃ�u���)��[�����v��gԋ�6rN\@��J�T6&D�ͬ�X>�8������hPV����u:%%#����=��|S�?t��UL��l�H�4e�;����H��)� �3���(�)���Q�N�i&L����v����t$*]N�.�����eB?�}.5A�*9��e��m^�KCo���C�E��f��J���s\Ȟ��6f�Xr�Pv�/{7i�x9�������P��?!y�0��B���d ;^Q��N�g9)��1��A�.r�Lӗ�E]�I�W�wlj3ZI�.f&K�dg�'7�|�3�
j}� ��!v�	�ߖ��e�ێ2#_*�? !7��"�[\`�*Ap�혥�����̔ɺ�&����A�N��	 �]z�/ ��j��q�,Ɣ^�Jh^��oN�/ο���v�;��%fG�(��Ӟ0U�ua�B�vs�j��)��(����sIbpOj,�ɣ����xCg%�5~~�Ql��.�Uf��bK[v�x'�0#[�/>�ߟV5��-�h�I=�$�Mwa��\�iM�bU��V����h2��dGb4�����AG�u��C�Xl��{�gT[��q�Ā��гj���@�J`O�NwR9�p��Bg��?�I��Xo�"#���pnA�u��?��0���w!6n�@�ߺa6�-܅�腩B����'�a�8�	W�%㕧��{�M9���/Ħ�<EM �M.�������