��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȚ�``�+c>�%�o)�`-x� �3�ڬ��T�"��4�Or�&[���
��4��
Q��+iw���zI9�)��\ڌ���ߜ��W����(�f�^}D] M�SE+w]e�&�Y}v���}���+R��w� ��I���Xx��A��}��cE0ʊ��<�8�⠔������-�-޻{�Bˠ��"�9�?���
;;����@�m!�(�)B��j��IXd���
�o��k�,�3'�H�xK�o�� �w�ث1E 3���Ͽ�I�Q��A�;����m	W(�lj ��X鮨�ʓx�)F�[=�Q�#���׼���}��ds�;��jP���XCm].P�J���(�?0Xտ[k(FS6Ǐ�O���
��6�8�*$�d�=��	UKh���۟��v�}�P<�yS�� ����BD�$�b�94��{F���y���j�f��ޜY]��� ���h��j����6]��)�RT�����'^��8b7��HkT���S��D���5��n���p�NQ/��ŉ�e���!���D ��ԗ���TKg���E4�PGs����=JhZq�v��G�V5�����P�C�������V�N�ཆ�����nT�9�tM��6a�W�g�����d�䳒�`]���,4��<�T�Q�֗bP�2��t��S	���t2}����z�[�`V��������^=�*1�ؖ=�����ښ���V�|���O��%۱0��q����7Ep���Q;r��`8\t�25�0�F�O��s9[l�G�o'�MpIc�l �ݽQ�U.~�'��ZM(���,7Y���~�B�BA]���8jb1_�I�����b�D��a�y�g�ۆ���,����I�L��6H�2{�T�dz�W4��P3�S �d�h�x����^ ��*I��啟��m����fk7�(b��,�_ 'L7�1��U(ej�tuX{{".��
�������oi�wA���ź��r�,[�5��0��1�.N��6�2�%)�iuj�^�ē$��>����NdL龟�Y��OC��9B��U����~.7��Pt4WM��K}�u�D8x���*����w�f�|�m	�:�.w2:"g/�݉kָ�p�$�q7�"�~v�7��s˽�?<��;�b���-�i�U�/�p���9�H~�2ս�*�b���=���}����ug@n�/����xO�ǘ�@�"��L$5qn{C�m5����Dl���	T��_+����.��C-bge~!ݪA��ł%{��%@�:��m��)ډ����}7�0��Bt3�*����R�!3(5��-�Շ1J��.�\o~��(D)�
��h^z�+��"�2|ռ~�ሧB��4T#� �	��Ż�_�9Eԃ#U�aW' )���<�d)4�̯��ϕ�a
H5۞�����r�,�0'��W�Z���+E���P�p��M��.p��}"�iy��a������'.��iP�#������6� /9{u�L�=�|m��]��`�6�R��>x7T�(��פ��I�"|C��U�Iu�.�iES�y�	v¨��q��Z��VC���S�h�*��[O�N�����>�N�c��b�I����h��>y4� ��߭�H&,=Ѝ�Ư���U��c���7���˟U��Դ�+̱���D��*|�U4h��D綟"��}�E\ώ1ߕI
�����d�bR�2�Je@ڌ�Q-[�р�^�\��zڠc־=?�Ł}����	�<��d�,�R�QW(]@�����ݫ��cz��T��!7��>��)��z������µYY���h]"�ɞ�~J�5bڶ�`�N7b�>:�=҂q��,�s��ޱeJ���3J襁2�G�͈�f/����9����%�f����R���`�`��ϭ1���TöuM��
^�~���vĻ�~�.��~,��e;ĥ�3����AE�����q_ (������]����p����M�Y^�f݅afdF��c��Z�o�����QZ�Tn�x��F��E��,떱aB�4��Ԫ}̵?�,w��D�RY��?�f�i��-���v��v���Z��ɪ`�>H��s�7�ET2$�jh)����#p�P^̍���ˊ�ۄ��]�_��H1�N�=M�!�Ȍ3<R����+k�ã��*ϐ����`I�̨�C}P2���Qp��n�$_��m)��)�\���.8���u�+���\Ѱ'm��H�?,e`���x.	�ֹ#B���U�w��E�r�7W��ѱ]ʑ���a���v�c_`蠶Qj���]�2��+o�T5�&⧓�Fl�r�H�>�׻�?���-d㖁.C�� �Q���}���2���N�n�)Y�(�$�5�'Z��XFw�p�ω	�����Q����f�eh���>�}�{
ޏ"~?:�`�!��Ӂx��I!a��[���K�|�uh��VX�E(sn��Y�φڃc�tE>N��&�e�وX�G?
��ɧ��(n �g$���x�� �"�Kԑx�&� Ӿ��v�X�	0�y���#֜��)�bU�ҳP�Bd���f��}��ښ��>�x�M5��p�0�"��Cq
��uM�QG�N��������F��"#�Iw�9����ra!�`�$Ȧ���`�Ǧ9DO�7�>�bA�̽OCp�zJ�2�]y2=���0J�Z���f	�E���j������yc{��F���X�?�w�c�����#���$g��ɋ�?V���7MW� Nt�h��agc���4�%;�>���]B�p��H�׻:D���7R3���1�����}?|�� ������#�]�~4��Y�o���O�˄���rs���ㄜ��Aܨ-R���+YK p���X�>�P$G*��ܧ�Ԉ�Ȁ��a��(����R��������M���#ߠ����YbП3u��o�n�Xp�U�y��*����E[�+l���9���$�4���Vˁ0��n���ic��=���h� �_M�Ig�n���\!/�H_۾\q�-7���%iNlaa)�E��!h���9^��/A�U���ްB<WA�nU2,;�w�2���_͍gG�3������������lp���_����c�xY�=�"��>5�/���#c����*�\o|[��Z��A���Z~f�Ң��W?�e�Ř��HB���)� p�fӇ�94��垍��i^��sJ�V\	���-bd,�O�Ǻ�Hs��V�X*���6�BF�'m���`�7y�ɲLt�sIY�ĥ��V�~^;��D����ѵ��ɳ1��&�9P�?m�8�#�ya��4��{���]���l��$�Wf���3RI����#����.SW�w�%��P�s2n��A%�$Ԏ��؊�x4�� �-h���}�;�`��p�?��?��#�V�^_� �M#vA���_+;x�~
��+6mKc�>56[�j���Q�0����x���O/��P���)��u�1#��}�y$Q����7���GQ:Ac����=���b1x[�d�5'�}�)�]s��T�J��G4��]X
�� 6�9�T2 Ȃ�x�p�:�nT��d��f�U��$a�� Xc������>$�����&�DB��-l2���x���ۣ�L�=Zi��F
��qW���R��=�����B��C�� �y�f�M���j��1��?�Eu|����׸�e.;���O�ŉf�Z~6�+գ+���YiαX�Л��MMW������e'C����槾���~�M2a'G�!P���n�O[��#�L�X�� 7.�A�M��dX��������� ��`����Z�ZF+�G˦-��,�.H ģ�B5�?b^�)�=��a�	��� ��F�r��o���I���)χ'���&�L���dCT%�sK�O
���,��vv��-����Y���8R�0en���?.5wG��o(PB��o(c��KÍ�O��w�z��gB� ���ۉ����H03(8f��^�X�s\<����ߕ2P�)�[`�[��k#b#�TP�+l{o_����d�ѵy\}� o�YI�ĥ�x ���b�^�N��oA�����Z�G��՗�@�����?.`��@Y��&SH��JƏz��C����R%�1="hޛ��Į�>M��|��=��)mk�r}N��Bͣ�y
���Ȁ�-�[Q�сw�d��3��F�,+6;h�A+�y�f/����@�+,֒An{QM�����Y1�!���������7�Dy�#{�1�V4ˮ�˞���f	�nL:����:��r��E�N��^�����<$���$��EC����Dx���AD�����Ӕ0曌D�V[;)4��!���/Kn�2��-Í>�W#��u��i܀�ǽā��H�}HӠ\R�� �E�:Y�	�9�
�C��&ǹ��p@cS���5+�&t'Q�9��ʇ#�1p����@ο�N�N�B@:�%XO�^h:�]%X]���i&��Xĵ|�{̈́�vc����;���v�]��j���,~�n��{S�I:����!ni��
M�Nz�F����7�Q{<�E��?S[�C���

��hכ�t�a�e?� 6��]}-�YS��D��
�K$�?��m�~�1��z�q��h���.�sCq|��/���N�,���|~ňY-���B+��d';��e����%JR#SW^���?p��� ��������@)�ʐ��A��y�1zدeF��5��&����<�וsɡ�f}��ø�˘���#�Da.�7���7E��t�B�tЗW7)!��L�A�"�f(�I���b����b��X|�� S�O�6�Ͽa��ɩ��[#���ցĀ��~�+��FݼV��=#32%
��i�PnW'{�Y+����1�Ŕ,�&[�4�vU���#�m���
���Y��v|;����=��9���>l�Q�~K��O��2�R�
��b
��B�0Sϓ<���sο����YW@��k��**S��)�=|�T���k�t����8�L�yw���A]��kg#P��է���D�0eʿ�8�ߑ&�p�-�~��r�«�}"a.��C��-�̃mT�y�t����z{DN���8D����28T��ѡp����[ٖ$VJmٟ��-ﴞ>]��J��d�;2ҬT*訓���3/ݠ����)����YQ��H)뙪.�[J�(	q�kLLӰ�_�!�^�	�-Ε��o��2c@�|#s,io�BP>��7Q��������ө�x�왓v0���N���)���>�͑%	���_鷀������i�B-^S�o� ���r?-B�m��>G��v��v�V�'c��):�n6k� ���3�ȣ|3�.6!�)=�2���g[���#��ǩn8��A�^��G������O
���9�p�@�	���/��@x�*���z��d����1#����)�Uz�4�Ú���>�{�x�r��$R~E��;����+�:�޵���n;��?�	���� ��d$X�����W��T�B4c���ߓY4wD�d��je2Y���nI"����)�ꖪ��C<���������i��fH���s�ru���h2�b�Z�!�毴k����;�\I�'�iξ��X�:�  ��������mL�@�E9x��ٙO�E;G���6;�V���>V�<'#�j+�Rpmi9 G�eۂO\5e��:�lZ�/�{b9����L>���g�#zq	�&����(#�����FSQ��)���ט��}ę�˖"2Y��_��1Ӯ$��)�q�n��C���i���d

j�V=���X�p����:xn���,���E�H���G�Iޡ~
�Ka>o��h�EM����j �`+�T�Vzlg춵�h��lJ��A"b��q��[w�4kO*�-�$ �@��X��`E�ܞ�tlk� �Z�[:����&�eܠ}�������ZX���asw�;G�ˆ��6�[/��Q�Co���R���C;��l���'��]m�����ZՊ1��O-x�ɂzU�|̹N�����P��XLH���u�̃JL��^��1���]���ć����l�8��6=�ΙL��L!�TҦ�@l�II)���t�� H�8�w=�W:�a,zu4)���Z~�M7�tÙ��d?�đ�L��Q8+#o�;?>�%sMP�I����2uK�s=A�QQ���/h"dðe��q�!;�L�C�N�N�K	�
���y�\�)���(���ǢT�,ʈ?��+`��L��A���m���BOHx�-�L��Q�8���7�[>�S�V g��̵���U��sk|�Ȑ��uȯ�����.�p��JF��9�/�0�������Fp�S�7�C��ckƟ��n�tX��X6��.�.��! ��'���f���at����O�b�F��ltP�!p߉���h�Y	h��k���G@��C�(̪��ԛ�M5�G�(�#Ev1������rr�!Z��j��>�z�T�몛��m r�&�I��^sPDuT�9x?>�,�(�58���28�ߑoQ!%�G�����)��7�
��ޖ�'l����)�~��%��4)���n.��������ZG��mֻ�F7�X�TQg[��߻�"����d�˳��M�����'o4������D��g_��KD:�!6�'c�b@�x��杽t9��+�p�{H�-�b�k5җ�vZ6�(��x"Z���*�H��W'e�J�M19�ĸ��L�!�Blн�p��y[+bn�m-(�yw\��m�<����Dr,�ۋ�����#8`��j����Fh�z�؟ `�'@bQ9Ĵ	;ƆXW����'���EJ�y�nF5���mr��$oV��v��o<Oԃ�E�ق��Up��;�e����#�*�0��;�xR6� ;��|��L�e��Y���k~Q���tgөT�8�����=�9޸n_��D��Fb�����v������g�Uj#���o4��n��7��e�8�W��[���!�����jZ+�2�B���̣���Cē`
!D�51�v�8�y���]�ȣ��*���B@e�3�+�o�������pf?��q�;C���B��rP�W	8�����S�jF�b��=�%��9˟\{,��n�@�7D�2C��k��a�8�2�@�W�}sgP&��)��ð�:Y[#`H���K$l�\�f�?8��@�}V1P #���,�B{�P�Ӕs��)�\�3N[H,h�B��*����𢸿��������?�1�y:%	k%�il*Y��8/��1e>L0��&�9�0K��|"�����%�\bʑJ���]��3�=Y-"��ĒL�U�z����r���:��)�_�s�~�_�ο��z#8T]���D��
c�Zc��*�d<����
��)�sH|)~_RQ-�:
�L�gm�����A`�QӢ]Ce�����/��t��I��R�F�	�YQ�Z~����	b�vC�fg|�i���,�^k���A	�x*�Z��#� �al(g����kq��
	}J,���g��>Ζ�S�[͐sCv��p+or0cgv �G�Fܰ%HA�_a�a�n��������'O���(�/-�.N~&(]J�����qn2�o�S;SB��%�;��<b���zC�s�Y���������	X`	ì���G�a�*a�UxA㕒����i"ݙ-a��"qN��c#�w��K*��lHN:����U��{ȭ����V*C%S`��z���84��m�|�u̸���ĸ��|ДCQ����A��{�N�.*�"r1R�dP�mZs���K�n�qі|�`�c�2�U�'\���>���fѱԳ��k�%=>�f �_$	���Y�nK�Cn˥��)� u��C�TIM��8�	�G=��9ʧMY����@�6S��)&��s��@jR��Hh�ܸ�oN�z��|�+Ό��t������>%���;��4��?v"L������I'J�������񔠄����3b|x��Z^��ܵ��Z����7|�9{?H���'5n^�p
��ep�n��덅�PLG�Uyo2:�^h��)�;�=�5����������	��\�/"�]�o�rķ�<�s'N��f}�v�n޹�b1����]I'�j?���Dxiհ`ӡ��
��!zi���嵸�~�\��j�x�]����J-�!���5�<�/l�x����2��t?�ZI/�W�S�=SRX ���� #�c��Y�;B[�v�m���d��6�۟z�,$Q+\R�B�'�Y`�>��S��HU�߾�^���Z�9z?L�y��::�s{�����f�����i���A�"��=/-�����2'lr��7 �􇫯�/�Oqh�]$	���Ѻu��6�ާ�w��W�@Q�2R�\&��)wk�\����O���Lv����7�1�L3"���I4m�sX��Pﭴc��?C�|s���n��8�+�!�I��,�K��6��@(��1����@u��x������C����ؐ��H� ����U9Q�<��E҇0����o>)m#Bw����ӂ�x���d�dڮ�bK'�M��
�}��0�ˠ�����d�c������B�*��߯Ϡ�����M��4\i�����2�s dix����^���'ͮ����o�
��Y8�g��-���qͲ^@��&��-O����܈`x}�Q?�j�8ʕ ��E���"��񸭯ZVЮ������#m��WJݜs�MT��|j,�e�EL]3�z�����W��raX�z֚.�]q"�n�
�̾QU����#F�/�G6�h�gX.��x�	NO�f1�@,��'�k'�I�Įr(S9�b?�W!A�˖8���Ӣ6x�\ǩ6'�Gfi?�	\��+��ot�m����5Q<�ٴ�.o���&nI'��:�8�e[Kq�D7A��	�X�cǧ+$�K	=���kU��v4(��y�*�%������g(k�L��b��� ^y��!(�7�o�_^�=.Y����nOu�8�"��2��T���*7k��|�;�|
���O0W8�ߔ�X��"'U����5�bbEe34?�k������
p���@O	��qFb8�}�b�����B�:�E.T���Ǐs7��kj8M�1um��TL*|'hq{r�G������l�v�p��:N<ʰ�0���0}t���ӧ��ž��1C��X3A��YI��Cf�F�+����4W�|jWE�hh{^��E���hf��G�肳�'{�D����tS:�3��[N_�.��%:�&g�/k��WMaFl��la��Uơ�.~�̑��{�9�ȧP���N>�5Ђ%����x�cE���P5��]��M�����.�������^m	)af�®�"U�<�^�.CM�q_Wn3o�` ��>��h%a�P3]��1����ӧĂ|Qo��u���]%���]��fp��IA+���3��\<���I �q�����׹F?��Ƙ��s#��
�2G��E�C��e�q�od�$�IO�MC9]�LD�a)��ws\@X;6��Mm�f�xu�/4�M~~m�RJ�w�~��E*~S� ��l���
	?o�46_�_&�T���]5f>��ܖ��>G#p�a��BǄƓֱ���`�`��H#�.Y�ڹ#ėV�8(�T;J�)����.���;�qV-g�U=�@�I��e�厰�}&�)�~�b�a�m����&�H}�o[&w�_���2.�'*P�3��]�-|8�Tx��H�z�)q�4��J<�Na0�(�IѶCLٙ�L���y�TW��ӎ�
I��R�Lk?�����a�y���,�L�G�H��'�q ��{��Iw��)l6~�u�k������dM�8F\� | Н�q�2��7��2g��*Zd���R���W�>�4f�Wͱ�ؿ�k�t��|=�uݻ����ƻOS�o�P��Z���ɞ�
}��=v�4�����菑ۋ�!���;�'��6Ԝ�dk9�gůn�<����",���C����B�@��m���X��,+�����
���M:`4�����iW��CER����� ֻa$E�̐�'\�m��(��D�,�_m#)x�)XϠ�sH.]h�2��뉴���6����\��}D.������I~$r��`���Tl���n��3��L�0�H󹝯�"�j�4]h0��]Q�x S׀3ҫ��h��m��;IG~�k�L
Fk�T�U*����VmP�m��U��k�!!�@q���aF��������7�݆�]�ү'�LР��Gy2��Q�p͌[��{��7b� ���7a�����f�����*{�Ĥȑ��b6R�?�@d���~Y�Ǣ�.n�nr�T��Vt��K"��GZ?}���<�uQ���k���F�u 2�D��Pu�?/���@����`�я�aX޺ R���V���7)�+�fw.Rc�#��[o�Y�
F�T%��$��f��M@�N�Ԝ:h��&ѡ�_FXd#gos��P�� \/[��� ���)y�g���|�K�,�x�� ��Ya+�!o(��wp�l}��E����^a�����S���_Kpj[��т���y����dܮ=$�E���1��5D��( Y��������Rg�83�<��<.u&�!��gi:ɝ�ï,�]
�Fx�^�9� ����7�(�8���H��e�2��T�6�"6��z9�j[�sBpA(�2���"53;�I���11zg֢}x~	�F���+�\���m�k��GA�X�T�9g-D�e���|�����=�,�X�u<T�U��s�~�_����O����ͮ1�هx��#����tqT�
�D�t�*�9ڳ:X	D��,�ê����E0�2k�ԟ\�1�����@$X5�'�փn����_���d�9�]��B�2ݹz�a]�r�A
ߗ{�(}')"�4P	���/��3�����(��/B��\��7t5�L��$`��;Z&�ڽ�����{N0�p?���U����TBo�[���>M�����~�f'B!�]	~�@�s�j�M�.D��\�$��"	!������޼���/��
�W�����v
��q"?���~Z��V���xUs2s2���8O�DS���G!�����8/Q���W�lG	��_�R�$�/r�u���pN�v����dЙan�4qANWV~�H�8�y u�u-dL9��	N5�g��x��O��<�'"�x��h�a�zIxZ�%����e�9�d�{���dN3V���;��J�U}m��i�9aw���i?�&���QE�W2z��@�t+lћ��<.��O�����s��l��ybntS~�5>�
�-?z%q��9��[��[M�yKm�����a[gg��B�!�1+ T���;��I�Z����Hs��L_��p*o<i�OqdNXN�b{,/��@ |��-U�Z���*�rPx4歭�[c�����Yc�<>Q��(-3�d���<öA�,�w�#C�t�B�s��,�ײ����ѷ{m}��"�'�+/��S���"UO8LVP��T�ހ�!�K�:��t�� cta�@Y���$�%��C�Y*dn�4}=u�5�@��8r��ϸ�ڄ�>f��q��ªW7*.{hZ�+%D4�����<�/��`��>W�"�L�����W�����Wu��cÞZRp7_�����2��ֈ��c�(��٧7�~E%���
��́�8����1s��ݲ�ݙ�3l�<Q����y�Ș."���IN�eI�l��X����~����YO��;�m!�i�+>���gn��E�\ �+^6�M!ڻ�6��v�\:���r�0��c��>�d�S��s���Gk�*��Y��Aµ ��Zn���Y�"�iF�
���$b��/y��Z3��!";1�j+���Ux �є �6f����9��0� h�w x����ZySӽOW�0�6�U}��D
l�}/CU�	l~9�^��'\]#x\b�R�^��f\-�?���J�{���^V�Ǐ����li��B�ӆU�1�|��aRJ}1�6�{�ݓ��E!��8�*������	�"!���-h{�v�6��-�Uvu3#��)�M�R�][Vz�U�+$��ޙ��޺Pflj����h���s$��Wrf?�Z�<�,B��c���O��v9h�ُ1E�qR�b����w9��<9(��@��I�>�1������Kr�������8&�[_� ���5�����<�I_�~tT�&��CB$��^��'�x�Y��n~1��d����R���.��t�]�������i�-|5�0�|񷩇E7\�3�z4�'�(w���fm:~�t��Cu��'EC"IV(6m8{��F�vCy\�j�g�(Y����;9���7�(E"D�=���R�iFeTg���c~�y���5�\�o��Ƈ�C�
��Y�?=H&N�;9Xz�r�Ź��-��t�fVA�nH|o4�F&�m��9*��Z�w�6㾽
�:��0-#�y�2
���.�.yyx�8�?�(`��q�A�.(1�o�EcPf�,���y��B�9�R+p�C?�Zh!$co�Ӫ\�/�m���C�qgkO.�5.�2|E.�#M���O#E�Hys�8�+��n/a$��)��Q�Y��XӴx����>u� _=���Yt ��[�O ���sh�k�{W��̘¶���� �p���^sab�`ӷP~:EU�
���|��'����,ϵ.������L��B1RY��Y�KF�ItV�{�2f5y ����Q��cOީ�M��z읱�hr��o�,(N��^��2p��ao��ZZ0�s^N�ME%u��� g��TU����Ygn"O�i�UZݣB�d�.��j��
M�������U	�8!%'����oC7���jls\�Gvp�՝C�d	~�T�\�G��g1�W9@�\8��Y�u�ܕ#F�;�+&Ax�!�����`��I "�pB2�T��^��|��י���~Y?CL2����P��ц��bfQ��@&}.���B�(;���i�CR&PlaWJ��%�O��ºE�qKH�yF���˝4){F�?X����P����DmDxՄ���&�*-�#�ZJ>�A^��>�Jz"���A#�#�}ݑ��>+ú�fYb�d^���v�����c矋->١��V��#�@�t��R~�~���X����P�D�����^���VOB��Kdė�����|�.���'ڥ�����/?(��V�$'z���d)��G�G@�@C����Ϩ��[�*�Hj6G� �C4�F���r]�f��`��`�� �`��%ڸ$p)B��_&'!d�����
��foT+P~�7.;�W�[���O��-��!M���avK*I��/���A)���~��E#�s��AO�g�,���q ۦђ���ǡ�!+N���Ʋ����Z+l7�L��^��Oq�ˍ)���9���M��W�YKא�Jͫ����3��oX԰�	��̩�� yFx$��`+2ާ�c������Y��H�@�����X[kԖ�X�|ab9��g_~��#�8&���S�ubTSz��\h��@a����g�A��ޗ��-�2�J�[Pj{r'Ys"c������d�w��f�|�-r��M��w���H�i$*Ļ(�Yڥ�L���7��sN�է���������3)����^�$*
��5>w���t�h�����xc)���Li�<�F��ɂgi��I�ֿ��"&�� �cSBmw��u����f	U���P`5P��D�c����a$$2���ҏ�?Q0�c%�N0؆���:�T��ʄj?�ݢR9�D�bkw�S|w�3ooǩ4�t��
���}���F�7w�Nd��ۢ�6�8�)�C�K�]����
fu�A�(����;��{8���Iq@��hݟ5G���糪c�vX؞�2'��rہ�9���~'�w&�r�Z�҆��U��,�w�V"��2-���RY}DO������ƀfSw�˲��@�V���E�V0�里�-�t�S"Iq4]or�t�>��x��2^[���*ϧ���/ҽ�&z�x���XY�i9��d���w��<���)�*���|����}^��-�V�A��K�jf�3��/�U�p���x�pRV��#���q�n���L�ʪ�l���f@bI���@��b���:w���p�k~4�A�^.�^	m٩�K@)RۅCd��rE�%�ד�ɞφ���otg�\S�3J0)��"���6�������A���\6�:�Q���@eH��c�[�����Nń��d��m�$`%�v\-1���K��楺�{����x��6T���
�c=����)�����Kj�Ƣ��Í������52�6�n�.�v�4���a�	>8��3���6P�~cCJ�A<�@'_Q8��b�뭂�ײE��qV�!r��Ȟ�������E���J�Ԥ-��jK�Se�Cj#��1��6����ov�ˀ�ỗJ�J��kL�㗕�����8`6��R�1|��?�� yJ�ȼ����EP03wV}�LÖv9Z^�W�G�p��v)���[��V���KB��u��l��_���OL�����
Ʌե*)R�3TAl��o��Z��#oѣ!-�`�;N*��`���R��7�m}W~g�Y�~�5�G�Q��Fs}�����@�P{���9�e&���oX����'�u,zF0)Ms���hd�����>�$Z�i�U+I�M���#a�՟�"����ֿDO��I�p�7���3{�GL�w{��_�C��G�jj^��N��$��J���H`m�{ZC��dJ�~_��ފU��V��g��2��l��x> �<��W��.6<_��Ϟ"����TeD0��٤�$E�;<�R�WA���B��ǱJ��_еQA�kKx��B�F�vȡ���]遻��:�<2�_Oix���a�'�Mf�J������pw?v1ppW�tl�_�5��`C����|Vr)�7t �*�������V������6�������KX?�>i'�������Y���1]å����l�9�h�Y�F"W88*s �JI{+O*�uǣv��ӖƓ���6�B����̒ta62��/�q�B,��o�\|%�\ؔ\?2�F45���e��sV-���h`Y������aD����y.�b��Mi(TI^r�yՂ�Q�s���M��I��u��������g��J/C֨F�K�G ���ow}��J��^l�D�X�~�'�z����܍n��7�5���e��*2�l���\	0כA��o /��½�q�ĵ��G��l�����Ӌ?�^���r33��F!
������@ٌ?���AisG�� ���D]������E�c��L�����uAd�����?���q;��z  ��n��~�A*�*�px?���x�����|��<:m�D%M��2<�~������Ȁ��f�+c�D���ɂK}V�brsjvU�?n�������ԷP��PE.�ʍ�0$~9Y�چ�ɹIz��ys�|�C�X�O�!_R���I�8�����l,��:aکo��OE�$w����9�&����1ţ
�����#��9	�\�^I&��S�!b�[�,Y�t�\���Ȝ����@b��'�ٹ�0�C=R$&>` /E�B���Vؑ#��3r�n�BB!���+�bN._����k�biL�ۙ�X"��Ѓ�� I;52s��K�v?�-�w�������f�*Mw��;�[��?G��!��v�#���	M,xηu���ct�˷t����K�ku�
hA��jop1��Q�Mw���%�B!�g��;�T������S����ƽk��S���`NV$Д�?��T����?�K�n����q�31(�Y���>�@]Q������xC��Vl�P��.�`�ۄez���04g�}�7�n�rB�ݡ� g�Xu������}G�+!�y#��mQ���<���i8�ߝ�N�kD�}hj�@Z��N�ikOX)�H�5� %C�*+3���3#�՘�Z���ۉ���7>]��+7�S��l/%����# �Sˡ�#�j+��g���S�Be���]d�'*vD>*��p��@?|��M�U�}$/���L���A`K�$e�	+��}�l�*���*��1P/�'ք�d�^����L���YJ�_����{� �r�4.�z��xp�C䟧�noq���,�Rꂄ�>���po�&C�$|��@�Ϸ,�noS5Ɩ�/ �p���>#�V�%�ۓ��}>٭8+�^7�/i��iN����X�5w� ���Nrv��Ka�,�&��d/,��[���}8Fť) ��+h��M�fHJ��%Oׁ�_�p�@q�,D O[W��E�7W�'R�pS��C�_���Fu�[|���Ĳ���Y�N]��f��������P�u�M�J�~�.�^+ќ#������%Ə�
%(YūCi�p+����Y(6IK�Ft�Ѣw��q�9p�l]>��u���&��j� ��J��)r��Uk᱗/���Ej����B�o��F�� '|oK�󂶎��Ѕ���:��٦{N( �![̪��ҹ��o�����K��E��]�=�L��YˣZ+���E��
�~	m����ů�̴�73[[@{/!|-�8p�v$��?n�d��������b�������A!�U3e0���R�20��Ԭ���>_��٪i!���
h��婗#��&��W�I_C�.i��Ȣ�
�H����y�M��$�j<�g��;ћi}�mȞ����nT��N@���L{H��=ǩ���LT>��1�����މ/0j�A�B�\Ŵ�f�N�Gη>�V�ށ��q�Ƙ0O8�$K����MgS�	����B�I �#��ݸ'����>Խ��6e� l5@uA1Z�JKI(�-��j��d�A�h%\>��'U�[h�2Gf�̠�}�P�[�W�ʸ�FԮL�8�%}l�o���2�"���%8��QE�D$*��qG�
~R<N���G�F�!T7����w������-}��-	|�0����_���Z[�.e�n�'N���vB�D,W$y��a����{�o�����Rw���R���/��p��<U�V�����zڻ~�S�B�s}�vt�����p�Q���|�8�r�\��XCIQ����0<o�c6�=�G�hM���� ����y�CT{O���Ѽ~=�o'd� gV�Џ!�%���3��*�˪/'AG�����RC�H�T���rv��rd�y�|���Gf�D�tW��^��cz�vQ�^���-Le���p{M�$}x"�B{��P���屈[�6N��Ja���ac流f(}����ѷ ��x~�-O�o	��� �rf4L(��W���N0 ���2�D.������]"u\�'j��ߴ.$�}���,f��j���*:�>q  swĪ��g�'�ɮn9�v!5 $ԧ�L���9'��s����A�j�Tm�y�:R�i�T��vѺ��V��_@��-��=���vbZ�
v]�Ɣ����뗋�u�Af���o���j��Q`����nK�B����w[d$�/-%����mc�ⱓ�� 8	ŷ>P���D�ZW����P��]�=�Ȱp8�{�t�����P�����Y��:��ʈ&���^Ĩŧ�=��o�A¶�Aܝ5��'�*V��/!_� =��ֵ�w��Z[��S>�"�@�5�ڞ���6�У	l�T�e���6��hW�Z�kw;�q�������ֱ��k� A-jZ 0h�I'K���B}��c��\o��8�>��/�Ds%*1s(?j�.xj�p�U���O+M���WƔ���/��CQ��%�J���O�p��y����
_�[%	$�h4��ub�׽������5cs*5��%+����)p&`�i|�N���=��j�{:xۼm�q^�L��'��V��Ff�8�`���Lp��C�V�,�c!�⣏����]�~�Lde��.0�%n!���3��aЁ�2'�_g��K�}�a��d��q��Y�vN�f���˚��Z������@�;�o���g��Gǃ:a��l��:y���?T����d49t���*�x����5��F;��o�m�oq��]A����g�����T}�b�C�伐�A�jڧ�V��~�c�H���o!�:�z8�{(��O'�y��&��� r�~0U
獗�=DH/�834�WR�y�^"�U�3��ɱ��a}�01a���\c���8���_`/�P��(Y�45c5R�s7�ph�J��tB�-��[N=b�ZqY4F�����UL���|V�*������@2�§�[�����H������
�mZG������j�sGȳ`�E]RBp�|flɧ��%Ύ�w��Qah�O������ƍ8���Rd�z*F^R6P�!r_��Gz�f�χz�����(�~�xCQ�}��1�eV����o:���0��Ns�(�F��������]O�!%��i�՘iÎ�_,�-Q����s�V^�vo�&�;�<�M�T���U���N0|�(��g���;�N�3�R���UE��f\:d�P���,Le?ΎM�;%lXpi,��Y}q��@�$#Mo`pM<�RS�����}��i��Uj���}>��e�Na9�j#����)�!�(sY�-Q�\�j$�zBg��¤Q�o*�����^��g��9���������׾�+�K�"�P�����n��B<�B�i�pQ{q8��M������;�F/�4nڙk�1è=
q��;����H�;�Xn�!8,��Q��%x/�s�L�a�f�9��,]��+ݯ�O�jZ~��/R$����w�H&�;�EQpɫ�P��ݾM1'<@��;�ڋ@x��`鱦���v�:U�
nBL"�w�F�+�%�ų�MX��>�'�Յ7�$B����V�W�`�ߴ��-����c���-ujC'�(�)8&�?��c��=䁹��*�?���S�f��/�IR��D;�_q�g�y)h�ݖs��:(�u'l�/6�)-W�(ʶ�OOݞ��%�]+z&��}ӵ`�q9c���1v�L�}/�)���,F����9�y*d������d���̍ku��^�n��C�A�k����{Wh�z=���Z�B'ĝQ[_�q��
;Q[�.R�D.�'Pj�zuHc���H���d���8c��t��5�B+��b�t�	�Bn�2v�N�WG�� �����5��ZӪ�T�������\,}S���$&�,l�#�(�y�R_sd3���@��	X��*v��R��D���S��`���ER}��>�鷱�<�#�ޏ�o�2`B~AKB ��6��cl��5��H��r$n���h���v���RGڗ�N���T��lQ҂��%*��<"A�6T"����KI�}S����3��>�ѮܼS,b��j	� ~�Jz�ic��n�pA�
r�z��*FV�'�MU�vW%}��y�>����z�����쐃�ej>#%G�Ӯ@��mcS�95I��-哿�r! {1��푊�2 +ո�$�Q�#�<�'�i�p��_|CiEڲgV�C[���s��$!��HBI(�^)���WL2z�K �[)D꒞Ό:�u�0�ϱ��by���e�����,��7��=A��<�b|:��RΛ[@�_�d���<�qNZ3�	��n�0<���f�����K5\�p@NXlPd����l�@(f���Zt�p�>����m���R�!`�>�Rr���q���V�ڗ�bN�bz'm�kҰ�E4�'����b��� �٦�>�S����I��a�wE�u���,|C;N��7����Wb�ֱ|����{\�+	�b4�o8��A(S�MnT��%_5<vf���i��Ȍ�?^�v��*�q,�,��q�uD��J�쀦�˛g�իEV褐9�˦,{r�Ώ)���3�%vN����z*�q6���\K����hh����������`
����a�U��|�G$���5�����g���w2=R*�?��A�H.�K��؊�f;Vpi��3���v�J��M	��n�a��}�>���2����ύ��1���۷����L� �������� Mߖ�DЫx���;�Ԉ{�j�
ġ�f���$�����.�9�s8ٗF�+X=����S�Ӥ'f��1 �)"�~�|������#7˽��i:m�#�K5�KZw�dUux���+��*�׽�C�
.<����k�^-_OX��l�PDf�nQ�ʇ��2�`o�����$Y���9Y鯗VS���T�Kٝ�A��ԦTȂg��� ���$u{�q/�iy4ɗHN*�<�^���}����KVA֮uk|T�a&�B+5�H���c�A������虞�t7��>�u1�~������<A9� ��@n?H�e��W�ǁ0�ۊp���&Y���A[71JPo���3y=�Źv��5�@�\�RmZ�#�R�(����	gn;9�R^U&"h��P���D�b�U�_��F6l�(��h+c���k9�g!^��4�45�ҫ�.�f9���Ч��s�ִ}l����
fqt�0�RC��S��[���O�C,9[/A��9����_|�gr� �tUe�@$;q���jN���/�.�_�#�W�;4
O�����TJ�m���8�3zy;Z7��W�Y�|M�`��F`P!��)�E����o�Լ�<�_�iM�dJ�ݧ-jNމ���F�Au$�7ɣN���1�	�u��=3(�J$�����d�_b��QRۺ��]g�D���������!�8m��y^��ްܰ˒�AР���V<���;i��v�^X+D��4׺i�:��,��2P��9Wn�|A����}�y�ܪ*��z�Y�	s�+ۚ.25��^*���ưe������{f&�ĉ��K�J���Z4ݸh�tp7�Ÿ��
\vEQw5rB|o������cx,X%:��ۍ�d���/`��j��|E��KMd6l���/]��O�l�/���S~�4���n�؟\RlHE1���J����6�����#�e����`v[=���
^M�D/(% ���Y�D8ͅ9sbۄ���+�i�g�N�Ǝ��`�}Y�F������l5b��šMǯ�P/��Kiأ!c��4�mM����o�~��J|������ͼ�Gi�K1�c�.!*E�H�&2� R4 x2j���q�k���^�x�u0XE�m�f�t��H�Oc&D��cq���i����,��W�Q�z�S��_wj9aK\���e�W��py�G.p����S��w鯩�e��γ������@ۜ%$��b�S�SU�`~�VD��bir��������c�>ຬU��oI��]q��GI��8��W;HZy�t13/|��#�iR�^��b]�OG0�ug���'��1W&|/��k��O���Y�ٱ�6T�*�">ؔ~��B�"Z�
e�I��}�	"]6 �J�AU�ԩN���FB�?1��j����䊅IY=}ӼHg�;.`QAsk�5ЀK���^���׺��P#lJұ��V�p��5	bz4�*�	M�ݑR,�)N����b��I �q^t�4�=�%���T'0�c���&J0�(�V�T�K�Y���DR��J��[U�1)�-
T�c��@Z�uS.�HL̀k0R�����}�r� �@���7���}e���T˱l�����.T�R.E�LL~���|�}_�ޏ9DE��>Ө�b4� �d�����ę�v|��6��y�zh�����c]
�L��|�ǒ��uk��<�A��O$�2G0�;.¢��^bPE����QO�_�[җd���`���ztO�og��$����r�l ��Ƙ�X�,����cb�R�p�ۢ���,Jl�p8*�U3L|NY������Vy�RJ�`}a[����V`K�Θ}�;au�*ޠu۬��r�h|2�^iH@h}��������V��)������S���#��©�g 7p�I�<�~���&GyPA��'/�
��,G�;W��օPxT?����6~<j�-���������^ъ��mbk�[4W�;D��랽��VE��ݍr�/�ϡꏡr�oU�WU`�\c��Z��ڻ�¯��'�0���X=a��mEGLIg�?!"T'���Ÿ,�ě�)]�[G���Bwi	C[n6�G�������{�^�a��9�Ys�,g7c� �z$�r%���c6e�1&9J�m9*>��Q�Z}_�&��fT �槠Ml��}����>)����ڔ��G:����DO�6����73�ƣ�<{��?odU�9O�y��XR�U��Wq&{o��_����~���k��7���η�\,���MƼƌ*��є��"n��
��˄�/ʒ�V�	�Xy�ș&���6�cĪdC z��[/J��د��UF����{�R�N]�DC�\��=���9��03�WtNl#&ػ��f� {~�����*/NU&1�u �!�[Fި��Y�wo��ސvo*]Qb��y�w�X��� ��{<�)�F��^���=�9)w�?E'#)ڙ���)*q��|���"������8/���p�#���4�	���}�im�M%H�(�Ϡ_s7�d�'�#8����qޒ��e�ٝ��/�X�y������#!K���ۀ����΃��oŎ&��}H
{�	E���yɮ�w�Щa�U��`������i���"�g��������ژ�����D��N�_sam(l}f����������ك5�`�>����z�t���Їh�˼���`�6`�_�.�[�r���W.��ɑq���j�7;��HAI�:�A�֒�����O.=9�Jfs1�goB�9/p˱�oZ���rq�6����Pv��d�GI�a�&ĻK�P�߽-o�7L?�z����Dz��I?��������[�s��VC�v�3�,	O�@u[���N-
3C�M�:��ө��w�g8�'|--Z�a0~�Q�[$y�8߸�]�4��G��{1��*�r�΢˩0�J��8\L�����k:Ɉ��Ě�GUԂ �������s��1��*Y�{%�>�)��������] �n��r�����[�ǝg�&weR�q��i(:�=�;5���oDh�P�٣˻���l��vo/w��XT��M�w�5�v�=ճD�c��CEW��	٠���"˭Ͳ��F
C�F�K�W���;it�v�/$\<B�P��a;�D�C
l��|u��I���K�P3q�Y�4H�#e��}ۖX�a#IR?jh���4v@�н);��a_�6�(��
W9�d������|)������va� �Rh��R��%x��;�&�Ğ	�=�)~���9�I�N��� ���Ü����|����F�#�ů��S�@����x�ʙa�2
�j1g���������oA���s��n��%������Y����O�ԠP2��6�-���*�S�(}M���U��T�sD�C}M\A��v��k����t�ΰ��2�e���5������cV����Y�	'��x����i��,�f�)o߂cs���W��r=ņ� �˲EcWqCb��^6�j2pI�Ud@��.$��G�"��W!�~�x�O\-ע+�~�uoY�p�� ����
3��5_D�3�ըM�s؉&���Ԁ�.����ş�Q\���۵�� ����ϯt�ze�)�0���Ss)�]�ܧ�fZ�J�\me��B�JD]vd�&=�D/��?g=簲�7�!�Dj���
m9��b��(�6-el����6�W�����=Α�@��3ߌi�k}p�I��x^���G���f��g���a�Qyv`�L���#Q�"I�+�?_EBlEXS<nz�Y,.�ƕ�7V�SZ{����f"6P��̤�0kA4�����6�]���]2��7�\�ɗ�y��L�%U��r2�鉡F�
�**�����8�L4}:�t΃0��F�9u%O��P�]�o��\�/�9ؤ��o`�Qi屚��<�}@�;G�q^t��6�V:�\��CА��cj�ϭ/|]��&�F��\�����q���B�i[XY�}csV����a�"[�[U�}r��+�L�F��� ��Q�C� <iE�ۈ��g�����:=EJe��@���:f��G��ă��D��p�M��r�^�,[8�@�[x�*�d���d�}o�S=:p��@p�¤�m�Z�����#�w�ObIu�Ie�ӏ!���*���*�ٶł6��kɔ��f9u;�e}�9�� BX��S�B%�yˠc�$��5}��jx�	V�W0$��Ά��o�㔮�Y��ATZ��^�)����7�1'~h�n90��W� L�/��E]�����ȥ۫戏虔�䨵<�(�7V'ly��V���q�Cu�m�[��]zu��%H�Ah?�����D�y=���(J�$�e,���veO8G嗬�n6dˉ�Z�E��aE�tL���	c���?�	,���8 ��� :�4�2��r@\�g"$���b���]������_��Rۛ,��j�9�b$k2��4�螓n��2^�p9_�x%�N�#^;w��5�q���F���X�#�8ޛ�0e�I��H�^I�
%��K�ϻ���Ŕ�{ۃ;�f4��b�t�#��W;�G?��9p%mR�,7
���z2h(�M�'�^P2�
��p ���9��(6�So���Ӛ/�x0�β޳)@�S�44�lk�\{�;FC�H*�.}����M��ɂ����H���=�G��G�Y����I[��ΐ+��h���e&�$e�c�3��q�~7�j�/�$�A�1��πPDX/�w!��O<��Dԙ5�3_�f�{n��4,�%P"q��@)hsD�n��������V��+e����z]M)�)p���L�Y��v��k�*�a�t�k{�';��c�9C�-���zX�Ҕ2�n��C�(���ҭfۋ���9����{>`��HF^����.Y�ҳC�f�G�:�S(!���M��ҟ���`]1/'�\	ѹI(�l��R�Z��F�n=!�N@��^Y�pm�UB�
,B�O!^=�ǻf���� ����l���'����+��f�g%2�}�ЬP>p���I������F+�/,�ikv%d�}9���4����r7&F�h�b��L�X˪r�e=}�{�pE���'V��}��x��Ga%m����+����iF��$��X1)��lJ���)�볒+���٘N�s���ߪ��K�5�p�tϾV{rH�<�����f,⦙W �-��Yr���Ω�"X�B/�/cy(�S�LK��-c���k�i��o�x�y�)�3���L
�F�S9�U�ڶ��Sk<���n�He߶���o��Y]��x� Jz�ܗ� ,I��Q�;��*��VT[ᨻa]�'��N�����U�Ked�a&�D��Sd���l�A6�{|�g@�53?P~��wH��-{s���dH$)�i��1�КC$�����,�*&<u�is{�4s.�4�?���N�Ƕ
�ךl>H\��al�(��a���ych�r�ֶ�6�H�[��E��n�
��$Л�^�:�Uh_
�я��<�]6�O�}%�����o�+�
c�4�g�	�'�3������K��q�գ�e�l��U��x]���y[��m�J�ߦ��\
Z�oX�n����u�M ��9>҈
��=
eZ�//)A�+;�s��o%�}�������t���z�E�	��H�D3���A��:��TL�����E�������5xH݋;{�ev�&�`�E�|F��[=��B��&��9y��W�P�N�	/��[�܏�h�穿��:G������IRZ��,�"s��QT���{�e�,�[n�z'�����P�(����/9㴼BzVj���qI��%ŝ��w$�$%!ײ_V=|��P���ݱC�鶪B�����7�mF�Y��)�&��]sO�m`�<"d�;)��[�U��ԘwQM�������N1{ݗ4��/&��d��H���n@
�����6>�F=|��w�>���30Z1f�?�PKy�����t��բY�v=2ô���ݏVw`70�@|���#�/D�.XS�y2.-V�q��zol�(�`�i;^�ra!�10�fh�"�_���Q���7V�U�e��BF����k
�.��lQ��x@a�L��Y��|k��]�����MV{������Iq'Y;Λ��meI��'�C�Q�x�z�.'��(ɸ@����>"�̥��#���$�G�����n�tt���bn�R lp��!M�eJ��oHa�xN��N�j��c$��_��;i�=�ΊWl����&G
Ƨ(@���+�S�/�:M3��1���S��H;�B[��챆��6^p�P��"�T1(�vS�[0a��W�ΠO�\����8 �[A�R��/��r �U{/������=2��}6B	��R8_r�3̗�2���h0l����k��G'��($�����ͻ��!�>KI],c���ՙ�������;!r���.-0����:[{�U�H Sᜐ�R|�ͭ��Y��\R�a�W��&9M�wYg0\�
�*&��V--®ע=nՃ��*�	z����G�ɺ�Sm-��ٽ��Qb��ԿP�����S\��e]h� Gg�T�����`��/ヶ{��D��@�࡭C4�K�T��p��|)���G�G٧"f��K������6$��NV<�������*��H�qI���ӯ��Z�JW�Y�@�蚧ww|��ض(��+��EJ�&&L�Ƕ||vn�7�.w�� e9uU0�X�
I�g�S���㊿k&��xp�/�[qܙ��T�:�%�5M����s�Ǉ��>S䓈��=��Q{As�9��"	5�O}��:��Ȁ�/8���2Lb�|�p��6>������~6a�t��<����W�g�t /{�L�2�mL�Й�^����0?f5Ƣz��UKFV
OT��{Ғ��z3Cg�Y��	��/�={�Nn��*H7hz�܁G���E�;���v$��K0�_� ����߼�*�;����k�ô���ϗt�@�)�'�_�_����o�d��h��ƈ�|_�XQFz�c�7��oi]��:z�ܺ���-��ݏ�f��CtT��|:�H���􍃉Z�v�k�&��	���:˾L�D�������ʖ�1��5�2�0��E�e�i����vz���y�<ަ�]�pT���b�I�mh��]Y�%|�[�=ӵ'����S��=�ss����
��gՙU��i�,$DI=щ��X T��3^�ϧÃ�LI;}�?�\�Mxo�ٵ�RZkp�;]��T�+�k���R<�IA�C�Q�������4���}U�UR�n�� B!�+���r_gU��:�^�t��'��e�m����F��L�0}+H���370�u�-}������1@��]p���/W!'�e0ҙ��B�5���5���g̓���60t��gWz��:���Vd����J�Zv�R�)�wQ��u���jZR�:��R�����5�AR�ͨ+�t�5"�{!Vtbʎ�=ꑬ��U�p��/	"ؿ��^Ʀ�m� 	z�u�y"�4�o�$q�Up$����\�yc�W_S�Vc����p�R�����Vb����\c�jO�Z�f��A�d~)띓bno	_ѝ�f2�^E�Y�3�@1��H}$C�qWТn���� ��F�L/�kϘ"?'2!�X��|M;�Q����w$�,���yOS^UU�sjp��7}'�������!����XtP%��Ȉ�<r}t+�(?W<Za?n˨<�u�!�=�ֱF������8�$׶�?�
���Re�c�?��OF ��╳�`0p�s94s��׹==�uT{���<��Ƌ)$HI�r�~��#)��ʼ).���{��}�p��k_&�L�L��=�K��K^|�t;�d|��_�U�>,_�=D�T����|�t:���"XkoT^?�m��pymt�06?p��n�/��Z��[#bД^F������wHйT���ݺ[����7&$8n!���f�L�����6�[�� ����:УS���BS�\���Zs�'�4�l���2�:P�P]�mէ��W?U���:)���z�xO����%^[!g[���]tҚW嗯���g:ޒn�:�d"\N|Ƀ{��.�l!Yh�i�}�1ԛ%��3�:�㈯�y���������JLKm��_o���]O{���	�>(NEYANR ��[��!]j�e�1t�����:Y�t����:Q���*��C�Oy��UYO�����L\c�ף����^e9�A*&�a���8�	!>�`K]~�`��;�%����z�ڭ�q�b���Z�i�H��WRa�S�M�e�E��R��3!��e9v%�n3�,�(�褚Qb^Z�F�"�a�}ak?�S�!��,n�����"�~�R�QJN��p�և}	@P ���Q������x��)P�Z�e����5�Gc6#Y�ma��L~aQ>.xh�/���O��pv(B������lp�Uc��#�j�=�\�L-�:'x��~�U.	���r��N2��`�_��^_�Qvh�s �RN8����%�����cg�w	WG��B7�,��Hy��v>w��At/1E�U�~�Ś��,c��X"	,��ws�����W�~y�(����h�:���P!]~g��NN�bD�{���{�9$��5;�]Z�.�Ng���BR��G��}@'�2���=��'a��B�zS=],Z\؝5�/~����D�$�C�TD�̎��;J���Q��K��h�3��vUq
xoG8�/����Z�QZ��o>z�/�N� #*��I��l�Wq7?Gue��4d�E���&�,�.�݁��a��89%�*Z*��Cd�d��6�WF=o��kXvH	P~��d�-�F�s�kD����n�z#�5���ηt,{���9sVb����H�w�_es��x=�/��R4�Rd"E�N��P���z�$i�k�j�v�@��E���ǫK��퓍e�^Ksm�8��-���VO嘜;nE�ON�˻�*y/G(�o"��4�Qg'��!�ھY��{9j0�
k*aŁ`�C�чԼ@���,'ǚ����/�B���=����w���"��}�Wh�j�^l��8V4�8���ܓ�S���;����E؍;�v���?%6ql��� Mk҆��}����R9�;}^u���:CR��M�ᭇ�	1�~����G�����G������G�v;~�S�:�᳖9�*�3y]��Y�tX�+ܧN1.B��TuMk<�SJ���҇��RB�Ң	`UKS�ᡤ͙��Qu	(?�kM��>3P��Z��6.�Rp�[���y�[�/�>���~@Ɠ�%!(��ѡ#�&�k��� �g_i�j\��8���M*_*�̗F�bHn� 7�����[�Dfn�)Z�{t�{��_����#N>s���n ����j�ӎ�\��%�oQbɃ�U����+�
�R\.����"�7O�x8PX�
�Q������R�/\g���P`G'�''4rۅ�+c��ʲH� �2�]Ѻ �_�C=��f/�v��'�O#wȈ^1���- ���<)6���c�����,k�� �Wv���u�!���)���Nz�Kp��� L0Xa�����8?<�nˊ�j�PG�)�Gɝ�m�k�l&S�Zhť����K��NY�I� T�tA!�L��3(gB��Ԛ����p�K�Z��u�p˅�k��0Y�E��� ���vq�_)p���}vӓ�ק��J��򼖻�F��jW҄V�у�D��;a��w^�3����^�+�	5.�I�Am����J'��?�L0I���\�L��q*��E�s�cJW�KGO��Dʟ��1�;+�}�1/F:��j%��ǴWSz���|�4�'�*|���k������~��5��(CB��9I�ͼ �i�)g~��R�"7�V �Jr'=s��Db�A'O���M��SÅ|e�� ?�6�[ϔ��� �1���H���s���2���7Ir�a��M]Z�wٰ�����p8����	��{lVnO~�8~��̼�R�OJ����@=��K�SZ��9ν}�"���ӣ;�yS7��q�A��u-N�jE����QY���h����r�	�`�"�?�j�o�~��^v%
�a�ێe��g;�  �k�b��^�J��Z��"��w�d���c�K+�� �U.�xJ3,}H�Ǿ��Te���J�EJ��3 ����8��rNm�+�Vi^=�G��Ubs/��D::��}��-��W�	��Cl�p��K���N{G Iη�����pg[f�T|�٦+���u��Wm�Z�S������<KM;�{�c�̡��x e�����]�ۨƹ��t�&�ݕ�-�����S4��-��_և�Ǣ�SQG':?��M:���g��83�6�M}��Jr��=C���uv��QL���#k�i���w���"E.P�����,,p|G�~�Ch�����)Op�oC�	~���o#����^�)zVB�9e��g��W�2tB+vͯg@1gO'=_�%�o�g��Z��(���<١��V����	ݨ4��RxW�6�vA7	w�ٿȐ�e����f#e�xZ����L9�O3���Ș]��Y%���(���sz�*j�P���8�Pz!��v��Aǳ�%0wA��7k��6��A��@h��q�γ	��كBü����>E��W�]��� �9 �{?V�����1_贘�,!�ŻcQ  J���J�x!��N���$J�h��;R  �h>��0���՝�:�]/��y<s�2������T�V`����	Ȫ�S�)+i�t���rb�:	�ưiM���J U�̓���JM��R+f@�N�F\��j�7l��!����aV�3%������{z2��q�׸ک�1S9��#^��N��bDַ�3����5T^�O�N��6)Ьu����I�"&-��Dg��=���`↗d�I^�j-��2۪XȽ��x]�4^�-U��'&x�1�G↣��_+�{9*S���߰`t�zXQ�K�Jѵ��3�`�H�rY������ہM�{5��a0�Eg+n�;.+�oN_���m��l܎H�a��O�h%6��Ap超���ϣ�k*�Ү��̈́q�~ۘ�4�[�c-�?=�1n+܋n��*,�Rb�=B~��u�/�6���u���ϜQ��P�f�a�N6�]Բ��=���n[�$���x���`RjE�\�#������ү��Bj"�+��r�dv��i�����+s��x1�y��#������X�{.�2�����9p�pN$�~.�R����f��T�M���gkg�Qd�6����:(${�d�r�*��!��t^E`fo�b,>n���=��J]���k�G�Ń��6�5��\l��-������Y	t	2��r���
ybe����*" �W|�_��������x�rvL��4���B�DY���E�]����L�6�I�7߸���UF�������~ҧ���3����37��1S�h+C�	u��`rzM��I�=��u h�������i�����S!9t���@#�7�,�|�@|xZ�&�>������\gֆ�Bݹ
	ԛ2j赾^#s�l o�d�#�ޔA��~�׭he}L�nA(��^М	J�1s+�&��� Kƻ�u�;8ms�;�)}�����h+|���`���I&@�*7a>��ڄY�?�ۥ�����������bÉ��=�A�����l����:Rc�k�:w�^�?a#6p_���Õ�̣�o&T��@%��п�+��ݑ	���L��I���k[r�:Fg�,�o�gR&<ئa$F���?�Ұ&��{z��׸sBN�"ת��[h�� 6�'8ΙKp��W^�I�Qe��k���C��U	�T�nȜǤ��=@�?����tɣr��	k4_}n����G
��ƲG�9���f�/�s�]��G$�L0�x"��{�w*@����*�!g�ȇ��8�?	>X�����e5j�I�uH���<�^(��^L��r��`���kF8�����f�朗w:��$�T3t�}��q�h]��ere�^�엁%�������s�pp��XV���?Jdِqr���,�O�oʰ\ls�t�Gh��8
eY�cR?�kDk§غ�$��'��M���5�jk�����}B�:��ޣyf�T��&,��v����u:�U��p0F�:�_fQY���x�?��dr~�����N��k�1���1��nБ��ϸeMe�g�ŭ�,�jA$�r������j8�f;?��EuѼt�VnىNѪ#)}��]�XMj��V�_5OZ�Y�gH�r��4]k3�?Ҍ7����S+1�<�n�zKO)PsԟM�����2�D@�~|H1A�|5�J̸형Em`8�j�c\�?��{��{�jZ.j��
�WY��pxO1��E�6 $�_�~�Ea��|k��4]K-���l�T�tm
b[ؐ8������E .�R�-(��дE����μ�B6��;wz$�S;K� ��S0:?�eￍa�~��R����5x��r��K4]��梎(Jhdÿs����5ˌ;q�n����Qfo4�R�Gg��$hf���7�j�F��ޏ�[�pl�( ��!�gm�@|uw���������B���Pr�˻ųό��ű&�;�'s�Ir���'��@������(�N։��/Ja�#ۅ�6���X�Ч�|�U.��G���r��29N�Mc�--@�G��N����U��ۍF��9�F����G{n5��8&/$��!E%�M��#x�1U���T��B`8.��!�e S�1�h3����[�d��Kk���A|l���+���N�W��Z�hg�ʁ ?$H��$q�C�W�*S�Ɏ���\�({����dzeg���"�O{�,�(� ���5s�&U�vi�@�Ig�d�z]���4\M����9{�M�����+;'eaFELd\ExbY��cPO�����x�`"�MF߈/��&�P�u}��M�T�;2�3&tF?�D>b��lX�i���u�]	b�R�}֢�9�Q�������Ɂ�'�n@�W�`��6*���U���N��@i���Ľ��H��c'{E��
ߝDwP�.#����/��Q�"��#�pb���*�TR
u�,�d!Ǳv��#dW�u��yH�ù��<1Z*���S3^d��1�ez��k�"��ȠH��.����c���2�Q�v���m(+��nAϫ�!�YR��m��ab��;@LoS�.|m���+��1�����*�9� ���l�j���L�1��,���;�I�(��!wN��.13�2+�RU�F,�:tK�ɀ!U"_�����i9���,��,�9����X�
�r��_��o$��-d]b5�?]�&������$_V��?��:�v?��:�lh��#��j>���$D�,VL-�@1�����+�ʔ�ж���g��[~��0����-�^�q���C���Θ�I��7i�;B�y�3���	�:��7��CX�ܓ����T���ߖ_��?��mۘ��X��)�@Ly�0��,x�j��<���,Uo�����*�cC�zT~{qP{cf��H�g�S��z�*��@�$D��2y��n����#hX�i��Waz%#fC���I�Id�d�6���`q��t�!4���M��"
�Vs_��ȼ��o�FZ�(%~�4��ܙpT��)3=r�zD�k���4�Ǿw[L,^jի�"��L�c*���ӜP�p��[�&�?����$z�,/D�Gd���@��������7�
ed#�^-�\��)�;�0A���v
bҔ�hT �݅��^Č%��w�����O�Dwq=�w����0o� ��$����"@\� ���t����D�����
����QI����b��Y{�����V��Ӷ�#���>n>�L;��ӱ!$c�U�P˓�D@�N-�\3�T�IG mi�`�z�༕S��އ� 2֫�Z���bG�9�L��\������@�l�*�h0������i���{�⃋�j�A��"ׯ�T�-_�»���'(CW[<����&��/a֟2{�VG�ɑ�e�)�v�&�K���L��4���EC3��'N=ۺn��f!w,!���N�(��:A���3#��!i��Y9	#E�K��IV1�'���db؜y�� RG�oR@p��sF�44��_��[3�S�6���xNt�Ǯ>�7u�V��{�ۜ\Z1L�kD%k������Q�k.���p?�x&gI<��zA��x�A��_�wQ;��`�[n�af~�ֈU�L�mޡ�%�Ba���
d��~���T��v������i�;m��=P��֠rG�j��,�A�|	y^?�O�!)'���OPs��~G3�ʅq׆ƢΙ?|��F�(��n,�Ӊ��1T�6_9M�Mvʑ1�pF#���Y-��}��@QG2���g��$S��m�����}�PȊ2���Z���lnceP��-A�Kz�6�i����M�<��)��(�ܼ�a+����ѭ�c�%,F������#-��,��1|����3k���k��P�]5��V����	l�������I��`���A�QQ��G�ri���t�qPȈ����1���b��T�g��O�D��^.��Y��x���U�,\p��z�ASTw��@��<z��
yr=��ׯ���R��B����I�!����m��
�z颊8oP �B0C�������3�+C
D�~ؓ*s�L��y`V9�H{�;���R����I%�Nl�x��vbl�hƎ����Y���T\}j�5�������1��^��9�2:Xg�Q��`���ja =RF�rV.�����J����܁9���}#t��<ڳL2�doKE!�Ir]߱SN� ��V���Yht��e�KOp�Q���n�r��?�|�Ng��{���Cva��S��+�6��TT�;�C\)��=�s$T�W��츫����7�8�2P�r�Xy�bq1�J��D�0��8��()�o݅��JD�I4J�q/M%��E�Ylh��:�����P�)p�tZQzAD�E��_@F�L�D_��Q�&����A���5�]��6��=����]~Lp��?�p�;5rj��[{ZT1>��?>A ΄�e�ϴ�8�3V�`Y��F^�,9A4>j&Ʉ�ln'1㵹�k��
���Y���nR�vN����+x0��e�,�LT@�MNt��"�p���`�1yGa$b�΂�]���͏^��	����]*OA0_1�UW��!���� p��Ϛ)��Č�Ӆ�7��U�����|k��_2�a���V�(�"�O_FK!R����\�
�W<m����7�r�t���؆`1�����Ky�G��t(׸"0��38���H)w�%�t�Mp\RHC��A�Buǵp�fB�`�}I�	�oJ�3"����ų�C�l@o�h_(D�4f?G0��|g�PX����+��0��R[��}�؁0���$ɱ\���Ű��eV��r�w�(w	^`1�v�#�"a\�λ;h�x>x4�Ln��I����r��>J��0�}}b�G��4�(�N�=�x�1�i���J�{ ^a��Ky����x�N�b����$XZ��12h�!D	�8p&�����M}Õz+�+���Gp���P7��fZ*a��n��L�+g�G(�O1Z1͂g��?FW�X�u��;<�=�ƷLɶ�'��H�%�b�$�q;/���I�{T3B�r�2Q�<�hJq�.�k�+�䭫\jʡ�tR�y/{%�&�~2�us�-1Xx�%�"`���K̭s����Q�fÙRs�;��A״����0Qq�n�+��e����(����;���@dt�V��@�&�4�)]�O��o���g������*�wnxmҥ�.[hO��b|�Pzޘ*�Y���e�G0�jr���f�>�\�V�񊙮��������,�~��(*SЩD!l\�lj�bܚ����puv�����R�)�U[\S5J��"��"�8�Ŵ���.�Pɡ�5��֩	����j����q���Oda�@1<%�L�X��r�XkP3�H�=��@�{�a�%0�ƴ]�#�G:������F�������`a�x̾͢_��# ��TKQ�~)?>*�'��ŵɑ�792w�y�[AK��#��8�#3�_���Z��K�u]йD�"�Y��H��\x� '<o�l�@������	ak�\�����G���i>܋�eNj��/�������������L[���0�#VR�lIo~9T���?���m�s|�q全s'FJ����"&���72>�WL�},�z�x%�o1�����Kc���n����S����q����4�p���?@g�+��͞/��9�����?�����QY��;��l�N+@��I���,�c��!H�OEu���#�% �����b��WVB{����ǑDwJl�wZp��P9w�G�xN}��G��n ��	�)�,�fI�dY5<�s,[yS@���G�f�=4��Λl
XA=w�zH�O�z�[�PJ�xϏ�s8y�iR�s�>C)x �q�2�f�F���֚�!��`��@!��K��KCX��ԉ�:�RV�`��P��G%�˱ǯ�@�5Yz/#}���H��6�OaB*����]J��vh��y�2k��m��>��G� ��)3[6o~-[C�جכ9���d��~D��������Hid�>$aU���L�%
\�i$ǯC��_���GKynp��`9�LR����� ���oj�JHzY]x���Q�5���}�U��U�����'��?V�}�����7���m2ŹgG0fTw,7�]fe.�t-g�X�����@v��|jl�E��I�K���1�3���0u�\�ϟ�_i��ѯ.2�&/���/c��޹o�
�XA�b��`ߤ��6�e�� Sڂ��д6�D9��C�up� �0�z2�udN�1���	}��۔����`�"����
�Iud9#9tW#��B�I2�-΄��a�)��E���NĐ.^�*8,���0��˧X>��yUPG�o�
��Ԃ��r%w��G��(Dl���]8�@�[7<�Ɗ�ׅ0W���/��\.L�JJ��N�����d���y��-�L(Ӕ� ��ṈD*?%��,ƋE]J�n��l�P[ɯX9t&�>\O�`:��ʂq�R���U��+D�9��7�B+��_�OV�dO����O���dk$o�* � WPJ��#Ӕ\0��Qfi���e�y܏�.�[�_*`�配B��@X���3�f����0_$��k��F	�-tK�2��j#c�I���]�!8�UM�_��?BA\YEL+�h2�ΓLop�(��򹑺с!
�_�;�a�	�:�n*U�#�\�~�/<����}���¥��
���t曁�cП4Z�Sg�~ �����s��!�MS��n���ʓ+������|�y"��xX	�>�̚|R'A�Ƶ�OA��ӓ>T	�&/s���*���Kr���[5q�_ū���BΗ՘���V�t]�X��<,�ͷ���6{&�g�^'�\������O.4u^X�Iw��I�ڥus�;{��m>�.���vS������L}����Z��	9���Y/�nI$n��bwm��BU�WG8eP���
����#�E��BB:8�W'!y�1�nC���V��1�X8�.���d�L�:e�y!��8$�@zv }.�%���z��N�|��A��w�.̓S)#'wDA\�t��e`�3T�����|���q��j@�!'�BJ.�)�	:��g�-	H�cqʭ�)��o5�ћ�k�h3�{O��Zd�����4c�3YHɵ�=2����~�y�������ׁ�/�I����
�4�?>���\[f����#�l�I!2���r`\�l��q�����k�#�cZO�~8�8o@ �}Ʌ���P�&���kW9�[�{YV2�Z,���D���jj��y��π:����K\"�W�r
�Q��X��C�N�l�7��Og:W.�W&/-?P��ÌZ�p�z�{W�K[��o�&gb����M�.0 �Zcʮ hmP�q��<��ʒh���'#��E	�"6t�n|�t�NX���/t��k&x`�� ��\�0O�EبM��fR+�m)V
���V׾�V����-��E���
	9�[�N}?�:WYÄ�dmT��(#?ĭ!���z�[�o_�2�!�s���žr�F��e��\\I����O�y��\H�!r&�:�4+����ʋ���z��y��Y�{3yK�l�%F�[�}�o������B��
�eى�=�1�u�HXt>�>A2�%�s`M����Ѩ�_�T�Pٸ�.Zh@5I�sg�H�K����k,�D��=19�a�pP)˱3�Xg��� x�/Z��������5����^Ĉa�?8h|��^��>d^3[�����'�2�q�W���C0+�hF��9��L(h#~i�7_F�Y�4�^�{J�F:fO�,���rC��y)�cѕ�G,k. �6G���a��b,8������	Tc��h��oYr2w�����5J0��>8zv������ցm�b�U�^�
ʆCYN`4W�������X�8[F��]3�-�#Ȃ�*��ջZ�n��%�K�w&�����9j1�c�l�v30XLߞ�) 2Q�$���G\��q�K�N-����V�W>E��u}U��jyY����@�/L%	7��MrJwC������jO�b��y@��Ͻ8@߼A\X
����V��F���sA��)͹��҆y�I�9u+��0�R�g��C���0��z�Kp��Y2�GN4d��d�u��j�mw�@�8He�k�'C&:�g#!�O���v�@n��Y�L^��E�{0�F�ȭ3�I�aŌW'����h�A�,0�N���5���ˑ���t�j�Q���GSM���a_f�-a�V���Kw���0��~���J��܈k�#���˺M�Io�3�$��?���D�
AkV���\�t�?/I�ZR���|��3�žCZ�6��F�v�Kf�ou�;���M���E¾A��L�l����Bn���n����6
��pHn�����z��H�.lM;=�ĨX��g�*C�����`L�s+j�����m�%�,8�����׋q��C|����Ad ��e{�*Ӛw��	}�6f��������g�����@��N\ys��k�V}@+�$�W���R�$���7 �E����3؄�N6P! �s���;�陑� R~RR���b��=��l�8�B:PW�hFTu�/ĎKYcA���r,0l�H����`���mS����q������jO��<��fB���6��k�P���0:(43A�h.8����ܞ��Ǆ���9���}��[bD��胠g^)��2RU�g,��<>WCR'��W�_�rZ���cV��18V�mD��缉�ߔ��8oȸ^�[�+�L�Tnp.�AiԔ}M�5��R�3iC0l� ]IaNeY�KN��6�w������B.����\�FL��q�I(�%��ɭчȨ�� �5fNF~��h6)Uon�"�V*��]��,�x�`e��)TEx8&�|��3Q��P�������9S]9���!K��ܪG�&=ݸ0п2�#K��̓jo7��ӭ�}�Uq��&��V�`�b�������p��T��wE𷇘 �#^�q	c�}1���D7��	�z)��C����o$0��Ū��Bз�}Qd7�<RD�v�&�[56!G�6vʷ�-��A�Q� ��v�0�i��bJY��7�dt|I���s��0҉^����B)���[�:5��O*��xިܑ�fDA͐ªR-7tв��5��Ŋ|�L%T+�#�"缾�c"���D�)L��m�e8�B{3ഷu�m/u7X��N��y!!�<�SE�������@�3�K��j�2a�7Ho2�ɇ�L )͉	��<��Lq�
`�<_�4���"��0]e���;Y+�-{I�����dAk3�o{wAr���^�|f�brz�Q����l�j켗����y$"�a�UI?�Cr?%�[�D}�G��(�$�6\������fcм.p��c���<m�,��zӶl{9FY�x{��xed�a ��Y<=h$�<J������A��\�<K'tЫ�o5��7Xz]���~ t��*��	f�s�{�s:���E��>�Q�mKnڱI����-S�f�p{����r|Zߤ/���p�fI�U�����M�{��c��<'t'�V�`�i�ԝ�%�u���YΕ[VxO�U�ۚEq��Fѱ��NFY?�/���M��w	Y�)��Kf{�C�[}�sIq��5g���}(�&�m��]+�CRI\x���N� �R��?��%ߘם�Xw~9�o�l3z?ZA4N�H�r߉Nw�E �w���hs��}��G����^��jW�pǗ�Gyk͑��9�p�2�7P�E%�M!mya���}|� u�E��隧)�@�Z���q�ٽbRQq�P~u�@
������������ ^�������>�=��Y�։�53.��jY��;i���^a��S4\�'^�ģ��E�#��x��mJ��������CUU��)&T��¾8D�t����N���(#T�͑�R����ē��C�"����\�u�i֊�K�