��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^�}����}��i�إ8�gO���:hMY�9���]� 6��+nM��9]��ኋ�/� K�M��F�#1V왮K(/w��w�Da�g{7O��*Q���I�\,(D��ߔ�A��BJ�y������	��,���H�Bf��e0���ａ�͙l��Q���>�(�-��委Lѧ������Imh�����L?͛z���(��t`m�i}���O�E�H���V)�?h�`��|�.O-D"��/tFy;\F���W!�j��<�A|#-�v��fz'i���~�}1&nsI��f��[��O�V��\�3>��.��F�.*�S�*�LK���Gpj�슺��O�7���p�&Ἔ��g�X��܉�(� 5�A��g��H��"�ʫYU��X��:�6�s������篇
=W;��w��&Mt������>(*��j�������Sb��ۅ���N}x&�\1zJn�Y/�8N�6]��;r{s�j�������\"(gg�cE���+�Jr��qYc۫���\��x+ei^m�
�
|(�A��l1�El}�Z���Y,?��V��v�T:�g�>��ʯL1�˼�5K?+#����I�!I�T�y��:�qlJ�УH������|��
�t��N�U�������X�6I���;�l�?����M�4��L�f�i��:��7��F$�����e�.53R�7�,n^㳭�zš�ϧ^�O�<��n�@�I&?7��SƆ��Ļ�q�`�P��}�VX7�m�Y;�E�\�7'�$)��m�MD��v������۫�vJM���;�'�{�pq�o_��ē�`��S�$εզ/T�,�QNI�:���$����մ\��o"�[�ײ܍n��\�|8�h��0Sw|��b��A��W���02[)���z���Ҡ*��{� n�o���R62>n�nN�����U�����|ؖ�&���5�]b�����k/�1��� ��N��ۀ\�q�{��[�h�9fC��w�l��I�"��(��F1�m���S���b�V�f��^��	Tu��8v�5����L��\3-	���Tl�6�Q�lk��1�&�y�{���u#l� �i�7O���;�v��$�W�u��Qc����_�>`i_��W�VwlS\Ȁ)5b�;d5xf�nT9�bVB��8���#Kp�$20R@��5b��I{�Wފ��K�Ԅ�a~�Xq_\�بƲW��%����W ��~
^�X��o����~��k���6��{;G9�(��������N8I ������L��/�S7�U��P������G�ߺB�Lْ��q��7�X�)O�Ȧ,�롌�F��h^(Q\��WA*q3��).��(�z�������`G��#���0� U�0�D�x3�[����(�]��Z^@���{I���>^�Pa�߬ƪ�{1I��YgV��>�j�5
y=U���b @�05��d{�rc�K���P�
)X�a��\<��V^xp���i��2ܳ�����(��|b5�Z���	�GZ	�xSΓ6b�h�����o�{(�xb�!w�\gia�t��fv��CC%neF�_&ك�������}�mvi����[wUsQ��=��s��Ȝv�y���-��"����ڙ1�D�Ö�4tS<�e������l����c���@-0j�K���e��vK����P�߯�a�Z�}�T<	�0iͫ�[ur��#�ï��<g\�7;�[_Җ{$+nΆ �i>�"���%W�_=��{V���Yp�1Gߒ�{˿\���]u*ݩA2H�Ȫ�@Q��m;��K��r�&_㈥�0:@�MOn�O�M�f���O��ا�Y��V���t~��R��G�@^ާTK�q�_m�fL��߳��%ěeJ���>���U{l]�#)��j�+�Vu���Q�G�!S��}+��(�)S+�o�l̓���D^SC�ܔ�d��5�T���w�� :�>^��Ő��-m��:Hv� �P�n���! �bT1��w���n;�(���`����:�Q�v�T�G�:2���ԡlA���`����x�+,��9�{��=�C'`YI��#��,��Q?c��qu�dN],PVU���8�|b����&_�`�H�x˟Fְ����C5"�zq7h����|]ê��s���+����!����#^��7��mƈ ǲ3n�8�p۩Wӭ��5�~H���fї���YU�r����Y�><�B@)�ـ����y�e׆E��e�G��U�:�;��������a|�UR)����E��{�R�BϷ?��j�;������{���[���u�c���f��"�.��H鼉w�y�Kn����$��	�Pw6�cRomA�0N�"R�i����`	:�;���F�4����kW�E��/u����2N�K57��߉3������|�P8BB�N}�OA�C�gE�y�4K�v0����[׃3���k�D2l���a��ީ;ű��'|�a�f:5�O�j㶞�|O��V?�JP&�?��w����ݲk�g:������%@�`��y�_tM�@�+d���u��ý��N��N�Z���J���U��V�������C9�dz{(�Xy��Nv��B�#G6��)돐y�n��zz��x̒E���d[��E�O�)!�:�� �;�3~�	��"�+1܅#��ۿ��O�1x�B���]����F|�=��E�������;1�m��e)�|wr��S����"�p�ΞE3��R�w'B\��"�h5{҆��܍z��R�Cbp���M4�BH�ȓӦ�l���Q��<n�D<�Rc��OdXQ���r��W$��?�^�R3��yk�5�"���N6�/��0�!0ޟy~V����%ʈ�]��c�������/ ��z���C�����?�v�	��-5q���t!J2ik�ɕq��"V�
�:�����O��o�J�� !�9�N����&!�h(>��mMg�͟�k��33�+<�5o�E�I-nL�b_X�A4F�.�R�Fݧ�A���#Tf�hZ,�@\�@/���n�І9���I]ZG��0�0}Tl�C�N`�y�8.�� ��=΃��&Y?ߑ�q�F�ؘPP�Q��$Y!�ک ��+G�^#u͏�<�X��tL`��睡x����ðTX���CW�:��J��S��_���"0�_C�D�	��
 ��X�3�Ww��1saC:�m�F�Ȟ����d�k��A��U%e�sD������F\�f���ah+�\����݄}a�Ԛwc	�F��M=H��P���sh�_�z�sD?��з(��L�Cz3�4�D����GA���N�
�M�1x}��x����;�������FO&�(����ga͑$���w{C	�%�!e��+��tc#d`�3���6�wT���g���g�
U�/M���B�����[���Rao:5�K٬�[��
��"���kr���t�*爯Y��c
/_'��U�VyW�??��OϞt�]#�(�%�.]h+ʩ�HU����}����o������PL�f�N� ��k�{����4^x�n����o+:UK��Nv�n=��/�N���j�{c;�/9�����_����n�<m3bBw�S�v��x�w�
0X�!Ԕ$���~8�z���5�%�v2�w���_�dW��,!U6:�]no8 i����q1_mP�������\r�@̰
�l�|QF�Ң[�⇰�5������1�lI"�j^�
�ܸϻ���F�|s�2�Y�%x��_=S5���:i��D�F�4����k�d�P��jҚ��f�.yo��g	��Jg�n^��©ǯ���ς�)s�^��l�8�XB�D)7� D��2^�6�@�}�FtJ�� �/?-�xV@�c�"�.w�HCf�h7��u */��i(��-T��b7�� p��l�r�"v7�^�h�J���p��t�*Wb`��3B��O��,Ys'�'K�ڝ]���m�^�X������MK��WX|��fG`z@�C�����V{vr����ݫ[Y�U�*�}b9+���ܟ��G� ��C����XnO)������Im���9���\�æ�s�X4�
S�cC�u�v�!TM�h� 
,�}(7�*����"��$>���/�$$h�e_�O�_�<��R�N�P��xz�	~���^⡲2�R��-I�- �����5��"��i��lGj���!x-���S��Kܚ��|�9a�l*���{�_���!���j��]�V��Kc ^��J�����a-~�q�Ɠ��{u�X���-�64kR%�����VBF�[��)T�+� a�j3�8�qlf��ԕ� .x��g�&�R>��,��T���} �ʺC�B�&p��i�F�.�143�4��cP��r-��"o-��]p�kS�v^�����n��\�����$r�u	� l��P:��a��'���1<ͽ�g��!�Ю$��(�P�����>�m*Ϭ%�:� �I��wd:�m�w��L
|�\�(5�VY8ף�]`긿 �Z3�W�2$�al�����<S��v���e��^� ����s|j
��Ԟz������]����l���Ѹ q�*��ҍ�T���#��ڞY	���ȑ�Sr�Ik�-o$3�V��ʧ�6Z�l.U_K[|��Q_���w���BzM������J�YC���l�C��DAJ�t�0g3:�B�$��A�8��^(�)V�9���8�����kR�g��W2Ve�â��*��:v��p(
a�ޚ���kե�Q���_T����.oV��/ϊO���-J�^�����K��N��U��ȼT�/�y�r�UccרYF����ަ�I ���e�X"�?�������<���R,"Q=*��O:G��1�^�	�R��7����Yi=��d�D�PX��I���q`>a9+�7�H��68�Q��Y#�`��$�#��H��d�A=-X�M�1j�(�/q������;F]��Y6���^�O��$�:+�����@wd3�e_KJ��y�����%&z kႈ��dLY)ƻ	D��\�e�y����50h@�V).QfG�%gMq
����Dټ�g|�q������x�(����U����$�EILO�z�,����.�M��5��/�T���1�[|M�`�����j����'�X��2�\c�B�gD�{,��"xY��P�0�4�z=ǭ!ag�]��#�*w�����E��Lm��G����Z���+�4ҡ[!G�볒�*�P;+�+~ �ۊ�lo6�$������b�&Y{��Z�������<c�Y��F�L^�SC¶�ۈ����=�n�e��g����K?��޹~/�_�	��d�ب�/hŇ�"^ɥ�dP�8�����)⢩H)�υl�´D����}���ޔ-+���٬+=�tA�fT��
�N�����:ʮ���2(��@ͪ{2�,�aS���c�e��e_�-�����Tf�0n�����'�h��]8����`j"5U$5ұSPF>��%H�}.��8��^^������E�O���e��i���i�2K��W����.'+Jg���P���'�kBM�T�=h�1X��z�%��TT;Ae����/�9H@L��K���<��rr�i_�z�e�U`?�
C�wv�ʙ]^���m�d��y�%U�1!N�*v��G%����>��
Z����f@Q��+�[f���x�����8v\Ȝ'��:EF)�����4%�`�l�A����i*�G�^��g�-��A��.sj���Di0�j3	��$�[
AN�zfǵc�.:J'"�A!l#�G?k�sZ�Փ]E��X����m+�tㆃ�v)��o��nK��jm���=5_�]0e�����Գ��0�4�2f<Եe��qncI?�|���:~��a�r
������%{�H�}�t���7d�x��|րEe:���0�����*'�˚0?�0�6���D:�w��v�*� (oT�q.�A��{ʮa7���e��R���i�2���z����Tj����*��Kl%���kB����U�$3b��##+���ap������^�O��8�GA��ު�ƫ��-m�����p/�f��ʅ�=����W�T����#l~Uh@�c�ua黪����!���˨��mS;�v[�ss��z:h�׵��d�~rw*2w����I���E�o���ڢ���M��[׍T�%�5����Қ+e�s�/����"������P�N5C0)�?T$���0RN�VC �Q��:�:}rm�lvI� ����C�(���pC1!�@�(�����B���\t�x�rx�v���ŮJ茮�����Q����\K�^��0Y=x��;�!Y�=cdѬ�4��tcQ�_��p<@�����Ҥr���V���׀�����@�,�q����GB��	��<ŋ�X++����%�Z��Ռ+����A�-�KP��D���g㏻��u��w1� �)��:�����"�;/�/y�������c� .Vfb��T�y�[õ ;@������W,'gU�Жc��H='?Bs6vb)홣��D��	^��X�YS۟j|��a���R&�<���N�7>�d�Qbj;IF���)��MY�$��g�psUQ�#�eI�U����N�+B���ÉX��ʠ�"t���	!$#r�]��-�f��U�nD��׵���(Zc-y� ��#���Tҳ�g�'�N7����M���?vu��^��K��jr�Ա��O��8μ�o�<sK8iu�;��x�)�.�l(	�e��)�AsYL�� �]�uK��E��Z�So�2f�5�	��>�a��(��v;:g�>q�T���F��$�k�Ӟ���%fAIYu���D$�{� a�\DH�M���z��=[��̯��G���*
�xj�����~�k$����V�Jрo��(�,p+�SHd~�����k��W��h��5O��>cs��%1�V�&���n��2[L�}���m5�=06�5�]_��J6��q�^�ʴ�X����l��P&�,pW�4�[,w7�7�fa���[�H�ry"I׍^��'��>z�x���� N�W�Zy��M�KemVB��4sIe���F�k�ԍ�D�#7�eTܔ�1A�d O�s~YA�!I �H �9SI�׬�S�x{�OV%��/�@$�R�_�^ȝ��7-�����xz �|�J(�7~���m����x�b
N:�pً0����Ah�������p����gq] �p��k��79'$P�5�y���-��d��w<����-q`��MA�e`ɯJ���	,���:��S�-���,�2�LK����V�)v���^Y��r�(�M��R=�H�O������"�t�/4��2�F��E�����waФ�-��;L�5��!���FNM�B�S��)�ہ�]h��D8��J�����^���_���(}o�G({���m*����ܕ���R���_�?¯35�x�
j[;d�^2�����+�9�Qnl�?���#�7�CQ�;dQ5�g� ���
9H����	YՆ<�c�"(3 tW�G>T^k���SiiW�}�|����I�?���3�h�68Dɻ?�Jk	��?oKrZ�qu�\��I�R�91T���� �9��E_���eYjU:	��KݬA T�voy�:T�v茯	r���6���KQi�1�}oGh��k�V�1V�ʩY�އʮ@۠����Yn3���
��W'��O0D�k���U��c��X��z(�������SJ�BI��h(KP� 藢8&�I>wa��Ez�c	�'���X��a����krU�{��r�8�A�ij�\Hn�&Ƒ6�=$�C�ARd�g7�d���Yh�/B��Y�G��P�Ts38@Ǖ�f8��� Twy:��<:���\�@��'#���vo�#�j�̱�^�"���̔��u/��D}-� Q�WE����TT%6�$�ZQ���!���-RZ��:u,��X�>��J�	�t���|��Q��BY�'k�t�/���r�B4�o}��/���#��	��H�4�W~�0Y,zlfI��(f=Dw�?J*��L����E�U����|uy�Nܹ��⿴�҉���ly)��M;�f'~o�P��}������!����lA�;����J����E�±�)�0����;��(f,��5C8 �}�w�)�"@��֍5~��4�xd��H_q�]+u�p�*�X0W���Zs�����g�D�����q���y"�*��O��0�����>n�sD�m;���Ғ8o��	#1��EqC�s�C�ԃ�x(/??��syB�g		R�\>�0�f2y�UKN�ʨ����_1_���W+[�q��p��&��[���kB��Z-8HG20�����zt��z�����ͷ�Y�����Ħ�U�`Go-��_��"�Z�{��j�N�n7�������X74�4��!q�/L^j�ᙯhG��h�R%��0�Gg�h<��ѿ����&�޺���|�U��=)��i�?BШp>�Gl�xZ�݋�����Ԕ�Qb9�������$��@Saɿ�]��@�<-M��P�<*wo�/�A!���X����ԧw:qsk��P�מ �/�&�,���]��My���Ř����.s$�ϴO���o�v٘����9�{rv�C�9��e��:�?�c�0T�c_۸�	cj�yl4��3B'HbA���VK��o���u )ݏ��U�%��V��JU�!׺?��ƱSۙ���b3���Es�6�ky������͆�fU��_��X�u��ŪI�����ž
.��$���gV�ʡx�QW# �]����ƚv��8���㩇M��S�z���@�� M����J�+��RL���3:�Cx߬9u�K9Q2�Xx�� e3��l�nZ�R����Ksw���w�A���!�2S����b�**^rm�Ғ�Al^�̇�-�����[e�l7�P�} ~ ��$���u&H�2>	k�4�J�R.�@g��\�:Y��'�U�"_q�M����1e�/#�MP��a��!�����~��eKӾ��z�ip_���B�v/l�̲g�_5ω�m�|��M�1i(E�R�W�C�+ [^(�PL����6�����[�=쯧�����؅u��O��l!��^E����y�Sp3�B��#0qb�3��[�ڌ��F�J�S��L5�e���[�1��y���*:A���\�Y�z ���"��$��a@����l��P�+�`�<C�1%�!rϬA�Qu<c[y���;�`���u,o�'[��� T_`�閒GY�Pz�����W�����Err�F�L�ؘ�G��x�B�P;ܒX��&��k��W������k�H���zYn�����0
m��fq4�rK~��s��W>�B�~Uo���9�l������9�A�)��n6�m����nMb)l�qB�p�������:�Ar�P�����5o<ȓ������L�B��<B�6A��XKT��'}QmX?�
����r�i�T�&���_������#N��;sƇ�`?���$6��y�"|ȶ��	��ar��"�qBקq~��O1U�ѱZ�N�T��������Ϻ���FuH`2����6z<�\l����� @�����:�:�Z�}�oI�t,�ܚ�7�\�]zn��{a,XV�=��S{�;�h�į:��#��3���,�E�p�w@�sz����7L[����6A��	�ʓD��R�Vt�#w���wrn�֗�h��O��1'��
 �BvDs����}�a�:�|�/��m�m�!d����g��p�Vk�.�s�f�~�
F�?Eyږ�O�k�4����;+ï�hä��8�$��	]X^�l�-��>�gQ��K��}t��0@q`��:v�� ����� �ٲ�^�O'i,�ު?�:��nlp5KM���V�}8F�7�ǞK�"��ѿ-.e�	��agwx"J��X����I�=��<0�p4�]��K�\+�8pJ�60g�)�ThhZ���iH���ݭ��Z��o����'��[�E��[ASK��C���:�~ ]��c�����AC�	uyޠ{6�Q5L�]��!�l[d�� C�΄ BU�ʳ���������d�eJ� ���KC�`�.T�UdU�q� 'Ȭ誧:*��D&zޫ����gb>���f���?w�Z[>�� ��U�
X�i��#k0e� Yǔf��3�F����_�T�y=��R�@MH9��s���0� ��}N0�W��M�`��Vמ|�d������!�x�o���8n]ݜ0���+�m1₭���8�^�����G�Uo��ѝ���bc�D�pǮʸ�G5px����a��ݧ�a�� ���C} �d�_��� ��r�ɊX)��.۟%ih�d�*���S��w�$'�sf���[��������!?��Du;4K�yw�k����m���X�"�-�%	H���D�n?	
_����㝃�h@]�5�%�wq>���da�uwL��]�)��ɉ�6�ܤߔxk��a}a>M�!n�����q\)/L� ���3@��&�?.Q�n���,��J��H�ɷ{R�C�p��5��a�W'��e��s��F�(�����'Ht�2��������O�[#s��/i��M|�Z�[�H��)����H���R (^�6Olz$W�v��"��R����F�F���2N��3-A������"&V��7���h���7<f�V&�����5�ĥ�c��Q�kc��f�+E�?�b�u��8�J J��	��B�d��K���oi�^B:P��u�h��fHU�� 2�*��T�_��U�y�����t�k2/�U���{d�4z5L������� �DÉ@�g/�|���`�"JG�v96����	��cm�"�:K��HO� �$�,E������ޯ�)}�H�`Dr߱L�B@Wsχ�D��6`����c�����+a��u�j2�o�����,���M�a9i�ޘ1��c]��H�+���Sr����9Z�GAw]n]H�������|Z�3��y�J4���(N7�P�U�̑j80)����0�)�1c�E`~6��SV����y���k�ߣ�	[���{!���1�,�ǑX8�_���"�������\j�c�W�ܫ>�AR����4�p�r@_���j�\��Tx"���h7T>���Mq�%>C����H�.��ʃ��'��_W�-��>����5��`z5���`^/��6J�g��m|@��x�~!���%k]����ܘӛ=�6%ӂ��^n�e�mS8l�X��I�D��t������2��!M��ߣ+���j��[�����C��;=�1�	���c���.���D�5��$]T��!�v���1�I�EdD$p/zH!h���
���6D����?�7o^��[?U8�Y��g^喴0dQ�U	��DO�L����[ :^��֯��2�7����̘ �����3�cR,�l�uI!�8[btX�K˱�ٵ�����\��G`�25��g����7$D����O�_�s���
�}R�{Hg`)p�O��{����®`"������F���$���r�;�U+7�������rs�o�� PC7��w�������]�� �k���61����HO'��C9yU�Lצmı�ey��{xsa���H���-c+p�,~�F0��(��yX;�������yE��i`�p �K����d-���%W���6KUe���<�� d�'0��ܒ�ϩ��%�ĝF[&�ÄB�~�m4����*���#�s_tF�+-�k���1p&ǁ�}I�qh��r�) �'��wF��X�Pog�{��� �mΚa��F�$cw#�-$ݻo_�O���]8� b��u:�K@#ݸ�x��^�aǒ���+�;�֭i�O��Ԣ���sL��t�}��߅_�ұ��kc�]_z$����	�j߮1�Rh���36����Ҳ���$JD	��H�U��A�Q�OG�O�p�S�i�$wf�F�S���h����,�7d��Hg�fC��)O�M�jߒ��L�i;Pz�u�;h�:�3�4�G�9
�&j'�1ٿ�T%q}E ՚�`h��w�(�y)��_l��g2�cD/��F���A�"I�{Uz$WkS�p������Uy�%&�E������m-��X�C�DT#d����%�S7C���Bʍ��)�ԉ�2��2V쇟��C�1�#�#�I���Aݨ�O����`�����cİ�F�/���e�A����̈́Ok��EH[���I:
��ƣw���U�5J���Wkc�*����LX�-q=/�}�3���J��y�(�H��kz�w;zL%#�ux����?���r�q�X��U�f���N��j$����7��f�Y�<Or:I���IT9��S�[}���&�\d>H��D��F������ܺGү��W�{f��",�4=n�ӣaTl1�o������c��F��;Y
[p34l}?>�}��2�6�i�=�; �qy%�έx/�Ok��߰�-S��\8:1!�N�j9��k�ٌ��A�o��� ����{��gW����@w%&zJٳCF//8�FM��W
�'�@����!�ِn��wJ�Fƌ����ۤ{��@2����
�f�Af�P�́1��,�6b��O_�w$�*�}���r&S���1 n����.��+�ebv97�]��-8�D$��#�(C�HH�''ɋ�H�h4��S�Un�d��H����c��uZ��m�rA7.�g3O����孿fm/��ej=����m�<v��=-�_���Q�usy�p2�>u���G��-��hRN��� ��8�^��<��{.Є��o���NI88�A��xjm�V�# ���A��/��ο���6�Q�kP�����o���N]���o��;bD��q�yi#�G9��Ɣ��x���s��e�a�@B�wj��=6Qjx�KM���M�<2����2���`��q��4�&;�Ȑ�9t�����IA�j�3)BS�0��RW�Y�3Y��ٟpIi�����.�?���	��'4�
|�߈:�����7>M�7�ئ}ٟ"��ɔaǴ�;f/};|a����T;�c�������1y�u���� �e�<џ�_/����*���U�F���b�A�s�?ŸS܁I���{��ZX�B�nnٮ=����4�?�����z�8��J{�O(i�[9���b���#*ů��h~�Q|�p�ʒ��a���I�pib�)���}�Rg�7n�_��#���/�E���F�el�ȩr��̓�PGM�w)p��Q]�m�w�Ǔ�����3{ƄݪѸ��݃�z|��/&\m\�Z��/���?��
$���g�&]�2�#E�� v>�e;���βh7h�/��[m����G� 3h�.GB��
�Otz���fȩ��};������02���t���9�Ҹ�̓]������w|�;�{��8fP�}p���I�������D����C!���A9ڤ@uk\b�fp�e���g>$s�5,��HbI��M{����}��������h{��5�S���A#@Z{�7ɓr�n�B�ڞ:,+�m�d"Q�Ǎ�Z9L�ρ��2�K]gL;e�U�ܲ�>���x[ ��c{�2�t)���m�V8?�UE��-�V����@�¶��[��v��2f1�:A;�Ċ����&!�PaD�P�jqiO�6c��s@?��('�tKG��+g�ϱƓ�n<Cz�NT�IR��lM�̕k�V�N��d4�t��k�"��'���XR�@V/�D�8�(<��������Z��;vg�pYt�C�h��, $8pAv�B6C\��5��g� �Ϸtg�ΐ"S�%�[_�R��ܥv�/-�P�!J#�Hy�*n��'Cku?X�@B�}˒��U��7�� �"p�^v$�����Ey^uL9�]����ƃ���)T���M��C�*9 ���F�ë�x5k`��Y(\��BWLӀVrK� �1�m���^�N�l�tD�	(0k���|� K:���u�qM�
��Q60��h\���3�,�'�L�K,��֟\��A�F��_>F�fs̋��mV��U⒅������%�/��r}�>d��֨�!dn^rTCh�@�z��j+9{R�jLHؔ��%w�--c�_�5�ٓ�"u?X�n��I��-Y��۳�Q�{�R��E�a�?�а:�y��(�1MU�"q�x?Hf�r��� h�-�ڼǦg?��_y
#p&�H�j\��R,��a�.)F/4FC�$����D��׈^�:��� _�H��SXO}��h�rw�땠�פt�D�z�X�j���N���;�^���J*��;���;z�f�xa�}gZ���"�kTo���u�G�?��Z�ZY̳�+@�眔bcj�PC-��[y�
i0^_,�]O4>}{?�BF���? B�'��VFx3���3ѓw����v��TD�/թ�Dʹ� ��n�������:A�R�������Bs���JY�1�)Ϛ[=��d4��"P5dP�����{��+q�g-�|�vT��f��<
*����06��S]%�O��L�+b�e��6���Q��]���N2��x@��B������j?|�����ig���AMI���!g�/!C幌�T@���f��9WL�u��>^1�6*��� b��E�Io��u�P[\��T��W����B�����Ŵ���&����5�K�E��{Ϟ������ծy<"<��Ո/J��ܠNN�hIE��B��
��!�AB[ fs5gz���|�ʸ���%+m`���s
w3�܍�݂ܳ �+/�K�O�Ok�q `��[;w��F�r�ݓ�t)-oKנ4 ���l.����Y1��p��~��A �� ܜ=�U�6�Z��6�"C�����߮JQEfk�ym���
��ոq`Ԇ����u�HZ`vvp��M�W��vi*+T��c�*���?bG"�w��+`�Un� 1�d:�N�v��䗼���9��6�����}Dtk�������Ɵ��y�����N�H�o/���[�R���UG�SR�bKh�W�GM���*�//��1��Ωr�K��4(�}����h�em��	V���FQ
��j�6���x���9�@��I�h0�Y��07�1�/.�����f��S r@��?I�u���e�����{��N>&�O�|V�&�=6��)���W��������fwz��o%�u�XO{�_�A�C�s�<Y]k�6�
#�hZ�������9_�ͽ��shH�ӸG*�9/�z�њO↕�]`�wC8^�q���s��7�!��SS�G8�Ѿ+$�O��u׻6R+m���ŏlq� Ef���lL�Q(!��1�-o1��J쯮��z��S�1X_��J��3���������w��:�ߺ*T�I����/��
'(`�׏^�#}��kӪ���9�&�/���j�^��YR�S��i|/|~u;�I��gWCu5�#�;I�ޠ1]OoWTT�W2����U��}kV��<}A;u3���~�}��F
�;��?4�3n͍�Y�}8��?�jÂ4��.���e�+�'$yܘ��˭��J�d��W�JRL�Ʋ�x3Z#�FۅT�#ɇbGQ2<��[ȋZ�l0��������Z}^�%�q@���\a�9�x�-�D���S��A]O�	�หQJ`�D�Ǆ�TrCf�U=�s[�ת&�3�p� 5v|Cv^Wu֞I����vԔ�(�7�<����>˻����r��Q-��Z��_�?Xj?㪁V&�b����XtVamR�9Q.h%3!�X���>�n�V��>�z�Q��3䵉�O�ќ��KVl��2"����iކ`>�/!�ņ�=c��^�.���ۊ�b��;%�p��t��5^�m�u.״������H����Q��-xSz��$����RI��&���x��_٬N:
�MuJ��dx<.�:t��$7�p�kL�;,[BDA��@�p���"R]�	G�j�`j�L#n�@��|0�.�͓?Q 5��B'lRV�Cml�&�]�v��h��S���,�-����?�k��C���s��i��%�L�����H�P���Yf|猊B�f{���?K}�4����wsi��P�dst�}F���5N�uyK�:��]��0�b�z�(T�t���6�6��ڞ�
�ٯ�h �[�lL���M���^h}(���M�e	����ź��7�d/�s�3�-�2�Y����k���Es:�E�b2T䗊���2u�B{e���&��
�����.Q���g8��ޜ�G�óXϥx�j��hɮ� ��d�(A�%q6��-����p��=��H�֑�D�%s�a�;�7Z�Y[�
���DC��>*��S��]\�o*̢�VD��U��q���]LQ��1�7��A,#����� ����H�lI�p!l߷5o�m�U��8+ȵ�8����NA��F�`��w9I�y�J;����ɘ�E�b7��{B�G���9&cef{��K�B��v{#I���݂*�����(	B��vE0�g=�j��{,La�DG�����yU����͋A�19l6����˙�(w<: 󼒡�-��ʾ���沉���ɗ��B�o��,���:��@nB{�Y̴��g;�w��4!�h0�⽡���0��Z2��_��H����2���� �?����Y�"��t����6L}N�pF�Aj����	.;	_�kl�w�8:2�Ə ���W3�p��F��.۪w�d3d �VҌ���_?j�c��f�f�x�μT��6t.�|��a���LAQP���E�u6���'VS�X�=��iZ5��Ɉbg����7L}3l���� 1�j���x��=a����x���Ѳ0Bj��T9]���M�x'�g���`V55\x+/P��s1��p�,�n�g�/��Sc��Ds�� [W�w��N�X�Fw�֞T�w��ƹ�����Iƣ������nqǋ�3>���Z��@{�!։����>�[�"�y8�Si�9�`5
�!���*�u�=�Ȝ~�m�6T�}կ��5SO�&A�Mq@D����E�b�R[�$��_��� ~U�}y�N6'���Q�s��5j���\fG��]"�n+�/l�AK�G���q)S�y��8�2����cYe^`���wD��l7ql���G�\��j�`�����)2�Z����r*R��S� wҶ�Jg�&�:$������)DF��&��/��g8�i�gp��\;_05�z;CX���\�ȎQ��2l�okg�8���k����&O\0;,%L�&8���˺w3���	J����򝍐��_rڧ�zx֟����ڔ�)mg��!��*�-.y��&^��}h����1��$~�8c�:-���ݦv8l=L���x�����<Kh��2	n��i}�]���q[H<�51?b+X�[F�	V�%}-O	8��8�<2;{�1p`BZ���,�ʵdǰ�U)�jeE�r�U����4^>��U´Ƣw��V�.��G�[L�W���~8%$���c0E
ThC�?������q��V ����]�љ�ЍљP6�g6����Hᩲ��F��ثW��	���$_W�
�E0�b��C���uϔ��;�IvT ��K�h�Sr!E۪��i^a" ��tT=0��׶<_,Hsc�G��4�uw&���^(l����#�"$1��h� ;�����
����\U��q�_�s����y���������C�y�&ϟ}��� �}�TE-��0��gL��N.�ޙ ��X�u�i]d�8�50"e;N5C��+��I��>@E{p[�2��р���V�^�����~��lq˘X�!:����0���n�����$�������͌�`-Gx�?��mP�N��'a{,�\�?�9yO�qa��?K?�����5�-'�I����V\��K�~KQ�u��B�����Æ9[u��$�G��8�1>VJ�܀��묓�V�b�;�^��O��x���z�g�?:�K���-W	��3�P�$�?�q�`\j���.��Ӊj�I}��ab�x��}=<v�T@5����F�q�G.�e���Y�����$�P���o�P�KI��K�l��,I���%4Jo��1�D��}��ѥ�s�6�UfU��>����Z�|�awo�Y��{�ly���89�� ��u�x �n�W���;��p��t�֪�3iL��af���pH�x���q�Ȍ���਑C,�(fl��k#���@�D��n|���>m'%�@phs�(�S���юJ2�r�5O�>���#���~��ڻ��x==��;JJEw���I(��'�O�s��$ĩWÁ�(-�+�
��;�Ҩ�������ͥ�yu'e�3�>�ٱ�7�@;Jr!N�sז'c���_5��{zC�҅��Xb��x���̡��>.�����u�̑b]���
Z�;�-��F�7���ׯ&c�t3G��:vX�4�(��Ʉ��S)�V���$��{����u�Nyw��kY�y�O�ec�K�_�E���(�RH~�VU����ʜ���@�{G���[��1���������ch^lZ�<�'PJj,�?L��f�:�B�7�q���֛>��d����BE_Z4�5]�;<���S�~�\gK��"����T(}���6[q(��B�������=����+Wy*3ѥ��p1�?נ�qrX+Ʃˢ0����<���̲�/K�.���F0ke��_�h��%bK�[녒*�:NR��6�2߯7_-�������iǃfG1�`[���.?�M4�r�r�}Z��,��w�-F�%��q�DW�(�΀SjN���J��܎2��q�zJ��<9R*��P�d�����H�٠&KDƗₜ����
���~�O �Pz�l�+�b�4�*L��|�C�\���o=��� c����+�ϓ�p>��]0����}vz����}�ņb:C��M��GF���֥FA**���-T����;�X�"��G�b`#)H�<4��- ;�vKe[�|�0I�l�]�)�gTA���`&#��+�O{I�����p�p��0iI�O�t�8�p[)���3�M�L��8f��m�YC�x���z]H�o<���|�[Z\_Z��m���uV�*Eկ��o��2�T��qv���m���p�'9�؉R2(?kz��8-��r'#��ȥ���'m�����j��R
��l�%���%~o������� [�R[�T�h��4�%���]��oa2��n��
�m��!m��N�]��M�ׂS�L =˅V�7Bmr�N4�͠\��:#R�A��2-� �N�1`��"�=G/EEߓr��/=~J�J���C��(��Ip��߰֎�f��d��/�>���}�S�"E���	~w��f�#I=2��j��@	�H]NR��F�ҕ)Q����Ƕo��)��ܗ���0m�}�ǆy��K����V���/�iru��$�u�C <P�]�� b4oy9)�ɨ�k���j�i/����������]�{��k>VJ�o.��Ղr8W��`>�|�o����9�T�ጣA,GΩ��5�}����k-�va�2�o��՟�io�+eeӗ��#eG�e���2������晥q���aN�D���?e&��cI�J���1�%�b�w�K������(�܂��oN^ʧT/ޅ^��[B�b�<�>UVEh=l��@G.��JdLu�O}�%-w�Tvx�Έ>g�d	�k,ܥ���g:��Ꝇ�"�H|�-����e�ǚ	����;1� M<fP��3u�&�����q唏��y���D�]�<uР�Ki�z���[:@�R�P�B`�g�1�U��B�{�V�<��iBH����8��Οv%�nnAk�����q8�Y;R� l���ʵ��]�هkh1�i4��+:a��j��S���<����`���5��i���P���~a<F���QK�]\Wg}�O8͒܋�c͚�N��5�Qֻ�C�5I|v�o�b�+erM�]�g%���&x�\�pu%P���Y���K����W�m�i,Q'�Í݀��'���2����~7�L۽JK�1ڳ���MAZ��/$ٚ0�f�H)@���	��ֵ�QȮ�/ͯt<�W,�յI8����@�E�1�$��p�"�_D��܄�_2�ȶ::X����ؚ�[�6�nf�P�������(.�`UO�* �lrQ�M
m�@��g��ٹ�v�S}Hm�/�{.@�xL����{ ƿ����Ԓ׷ױ��.s�ޱ�]�\lu�HG�jk��nP��.Q��T�l��9��AS��WB�o7��[�Ju}����2@_�Fi5a3;��� O��C8��Y�jQS�3$�5BFXEީ.M� ��w�c31]�|l=����6�V	�#�lX	+����PQ��ag�Co��5^��QmsLU��B$/��r;:t�w}�6/�vW�K��]����� LE'�[K��������P��c�y��q!��O�Яrf��EѡLaB��!Ŋ��{�L��e����~Y�w�l��H_��~��!�U�
1�����$�xv��[���5�?����u�fW�(�C����W>����4�l��v�7eu�͢2�j{M�l�ҿST�n�n�zw�%8MF[}��������4E�/qe�5�g��~;ã��KC^���X�[���#q�P;W�=������巃����R���{t��A���ɥ�Iz"���uV�Ykg����ͫ.��>*b�����x?�ێ��om�������Q���LF�� g��}�f��t;�A�N��70�m���\�_M[�e�Z��j��*4I/���)`=�k�C�Ȍ%��v�x`͎���TC��Q��n�쎛g��Hvdt�p~�=$����YC��M�4���b[1g�C�-��g�@�v��)�����呕��3�WY$X�|u�6�3��H>����qG��A���ߋ]��N�ě��fvZ�o���!_H|}�*���O�d�M�Y1KȚQ�FGU��rewg��cc���i�3���<�ka'u�d%�!U��K������)��+L���Ή�wKH�r��̓����t����9��s[t��������6퉖ț�v�[�}��_�.q�l��fS���fؓ�B�z�,���ZCl?v�<	�o���]�(�f���\��pS8g��i�o��׺�S����\�����������7���1Z�OY!UGÍ�J�7��!n'_O�W��+��>��E�6����!X�ŗ4u�@����?[�a�����Ijs3/�p�D
 �=�>f>8���>S�Q��#4պ(��|��j2<w�.��wh��-��JY�aC�`���B�_����(a��B����' Ë�GhmS�:x9cVo#$�{;.YU ��N!^�ImS�nBMr�{[��z�33��J(��42���J�k��Q��k�K��0���>���7��<��EB<̈́6H����_J�)��͸w���z�&����'�Gx��-�H��z�|6�b��7��B���� �y��02qS�8~Kv�<S���HP$�!"$�#����0�n8YO:��q�h=�un�ծz$��p�d�I�e|�:[�������ɂ�ܜ��ca�)����T�B���A����&P	���)c��&[T;��˖t	u����۳F#!T���B��"��-�r�W���l;<�uO�	��[D�q����"�Y��&~�)�R>Q�KC�.gl��_�<sEǤ(�g�6[
������5�
Ԙ`Ǧ�0��k��)����(k���X��JK^~,����x7O�\�{0�<"�-�Xު����g��u�Ʃ�=#&f�/hC��'|��\eghWu�)��A}��d�����.�G�M/�qT$�h�W*g)�,�8�h1�ڰ*F91k�:��X4��j"��Jg��ݭa.�\�ś��]�QB���'bK0�}�)�fX�j��jybR�G^�������+Z�E��K�=fO�3�.z�v n��{q>����2��S�"���1i;#����j�7K�Q9Ҳ�o��{UO�G6&$�
�i2w$�����2��0��3%��!���t���G���O���5��xZ����y�삛&RXK����O#ʅTo\N�H~>�b;_�,�+]G�k](h����h��w���
Z2�̍��ꮶΈ�n�]+�Πv�.t;�	�D�� ���.�0e��:T	0�E���;���O��3C*J� ����⥆u-��]��G��h��(km8���u��}��a:g���;����%|�r-#�� !(���B-�y��۸��ܕ(5Ӕ��U�b��9{�ɛ�4�f�d�Dw��Փ�j��_��c���{Mt�l�7a�� 8_%@>�|[N�H��t<d�o�g�a��7׎m@��T�4˼�GI�ؤ�?�8`ö��G2m-'.>"<o�J���*Ȁ��L�P"����L������4��� �jФ��+e�C8�)��&�(p���3J��p�8g��%BU�i��I,~댒��8h(�$N�aYp�E}:x��4&
�B��h����v�t]�.8uX����z@WC-��?�'Ih� ���dҔa1Gtc�Yv�yV����5H�pjY��u��(���:V�y7�u���X~����k������r��h�
�[3��E(�6R����a)k_,	�(����n7 �`-,Na`6������L,U��5O�F�;�О|�I%�aDڽR�V:���t�}�PjKieio�:�-�㞄0���z7
����w����2t���翇�ºB�5�p��/�h��:H����!�:ń���¥��ʜ9��@'�؂��RX�AqI�n<;L�R}�n����)OV�#��.z���VU��F�,�����*�S��S@��|��4l(��I�Zȧ�C��etȯb���gɽ��<�c�.����
k��Q�;�g���ol+ƀD@ٰ�@�]�|�t��4�1��1���l�R5A�A��Ǆֿ�n�D+C`�T�ߍߏ:�s��u�����\k�_9@N ��:���'�`k OpE�����v;���W�s��X_u)i�H x�2�x�>�b���\�� Ǡj�����a3\ ܽ��ʶ��.���KpGP����~��,����O���#�j9����ߜ{�"i���y����)ӊ����t���V�i��aWo�sd�+�?�wK�ѪR��]A� �7-�k���8�	[w�"�����j%v�nR�1�Yr�M����##ν�lE6Gu6� %��;�����%�}����踎���MB�������AR}�J�d����I��>{���K�?�;�P<;�{�O"�خǫ��{Bz1��[Yڬ���=�S��O��>�Q'{�&�(�l�|
�����9L�:
_z덭�?�WB�0����7�64�M����m'�g�����<���Źj1��"�Ғ	PW�0V��J�QO�R��n_wy��K1U��������?ls�1��#*��%�4u�Λ�T���w20��w�,F�f&F����γ�x�E����*�q���)�)n! 9�1Ml1�����	e��SY�SJ7Y�N�z�O��1N�>�K ��R<$�����k��o�&�xuh�ޠ@Bmp�������3+A��P�X�Y]���y��:z���f ��Ң����@-A��6�3|�Y��`��������sJ��ulÓ֩V�����`�Sc�����0���}O�D=mG��9���=_����dR�<��m�����?�RzH���	����7V�J�e#�c��P����ޒ�ֿ	X_���"D8{��5iF�|����T�{��U��o���KB����ޤ�f�<Á�n�&&���ȁZ�C��R������HA��ry���Ѿii��=�+s��8��	&G��䢞�5��R�� R�D
��8�!�WuL��d��j�&�#�~*���ys��W��'������~�4��^�tN�K��"M��[�BfI7���@Zp߿5�X(3��<pj�YI��	k��Z��~����ohسo�9����6��PH�(|ɑ��u�RY���@���-��а�'oI,[~�F��8]а��[숺��D�(%=�KBs�}̶3�M�T��a�X���&�טN�\�F3��&�k[L�[�����z�m�"�(��XS�C������
�졳�pn.���<�y��(Mw�X ]�f�M�U~1�z�@V�b���g��	�Mߚf��ϻ6��#T#�>�j��fY�ٯ�·2���VZ?{�:��`��	imɰmY����X�"*q���q\�j]����t�P*���'>����>Z0u`�6���{�Lbmw��M��B#����>|����	��m|��v���:�J�|���E��@.,h�+o��=7��p�T���a���n���K�s�I��u�	��'u~��i�������<��y8;f���[�o�õ�sn�b���p�u���a恈�Jz1�Ɔ���(&s{�}E�
�T��8���E&h��h�)2e7��x�7$����8��ELwy�z���WU���~��M���Pq���eG�t���t��,�~pt�צ(}6�� B"����]o�.Sۡs������J�1hbT	z�N%&VE����n�0���[�u�<_cD��ә�	���=!/U�Se�[�Z��Z�k�~4%Ќ��]c�������d�4���g�)��u���h$�|5���1T?�K�(�Nb�h����*�[묌�����8�\� ~�6L` ��
��pIy��'$+�3����U��<��L��-��q�H��,�(O"��ȫ�&��ǐ��}c����Q���5��^��h�է���� B�w��Ipq+/�����x��T���4��(f��}�/�s
�+)6ҋ�y��|C��ozQ�������β� a+��k�ҝ��i�z,(6|�2r���k��N�芿�Ԩ9v�.�\vx,p]˂�����j�Y�a~��������R
l��OW��<Bt�s�T8��	���\�5�Yg���>�]<
��DL�[� �P���W���n9��
�J�8�2��0�xӠ02��-ܒX�:����/�� �>�W����pTh.\	�fK�-a�y�!�������K<^L�ȃ��~�1��;�2vdQ�m�]�⨕um�Rr�n"{�"/��k^���.9'�5���QE����N>���� �&x�{�XL���#2�n|Q_�Fq̒
�����>�q7�m�=�{�����(8���,v�ڭ�l{�5�����Sy�~Ǜ+2_;�)eo5��uO����+�_ݱ�D���d& ���ʾ����l������4rM���?�̖|�������1;6�����7�݉pa��_�. '�v$�
�p
mҗ���`>��?M��y��q���t�o/���c�Me����dTB���&�?�IϹ#�l�/�K����F�v~e��*�K�+3�Z���iG�|`�G:Ζ[��g�}?�(_G,Ki���+n�($Ɠ�`b�ȮI�_�WО��5�6��:6
-{v� ��()\>�D��&\r(R��g?�)V�	�t�r�VtbR���;��,����2�ϋ!Xv��
K���t�%�T0��!R���*��Ng�M;GDݩ9ne�8"�� ����)i.$�&0�(YU�ǈs�:�p��rP�?�Hr�޵�6^��.5%��_k7zW����vp�y�^�<ݜ�%�o<��q!��&�&J�sh��z��Sn����l�V���H�b�m��}��R���P�V�h���Xzņlq2�9��J�זj�D;����-�
gH���S�']�Z�Ρ��m�F��1'@cQ��0�xvĂ]���﹥Hi��+
��f=*����I�.�ڡ�&!!��F�4��a�$������T
aiyL�;�� �D;}��͔W}�+�:��c��Tsʨ�}�E�7%B�~OJ̑�
�f	�+P����^��p0�pF��m�R0F��Hw�Y���t�ڏ_�)��R,VQ��@f9�� �Gi�|0�[#�5Ǜ6<%I�ـ	���m;Gi�މk�;O�)�D��,Y�6�Kci�xs�y���Di�_3�N:����3���[���%׻�y���"����.Rm��f~�^u4 �`"�E�d1�ԅ��qUV���,H�Z/x둚]/]����ký�nN��c�v�k�)�oj.h�`����I˼xmG@(�b�+e
�Y�d�ƙ���P�:�n+gա0�e��,b�2V
�X�f��r���M�o��޽�܈�.���
+f7�X�N�}��ٚ��l9}�%�M ��K��i�s� tӒpm,nN����Z� G^6����yj�OW�K5N��p�q�l#S�I��;��Yr�>7l��V����ѿW�����ħ�8V��͊&h*Ԑ�H*�|��{l(yD���d(���@�t�[��v�OTt�I7���f�1vBh��B����
�w��ڙս-Z7U�	�Z@�	�gꔨ%!�Q<_'�����9��?K�O��Z�[R��2mb�e�"��\�9��U�.��+�0��C����7�p
�w��L�{&�CA�Iq����7CL �U/o��`�[���A���b�'�|�	��	����8��6���ǆ���y��n2�W��_+0��&�U8�3�r����z����*����ܘ����g�o)[��p���W '�}����}�D%��D�Q����Rh��+�ط1�n7(���3E��BM�G�f�7'GEtK�S;X� )��ۧ*K�ibN�	�0Sգ�d
wR�6��$���t�O��
�����a��ۣ2�c�l� Dv-z�p`����kV�89Lh���z�?�?���3�^�P�{��|�ŝ��
�͒�c�[C~��t���n��\4ϒ���}|�ۗ.�_)Z*��M4OT�{B�y/��=ڜAdB�Q#�"|���y���L�op��a{��x�~.��"���F4�g:��e�p>�40�J�i�:T��A:z�`�9���]p�(��s�=҇�R��g1�Z��!q��� o���ߙP!f-FHA�Dԋ���Ϛ�� �"Z�|4>����:�O!� ����Ȩ ����#��3JB��pD�So\�BB��g��7���o ���I�Ƥݥ-Io5�1�)?��T��$'�sD��!f^�}uKOo�৬e��������'����Z���Ѩ�^]�m�:,��u�����4:����IC��bS�!�6E�����l���u�9xDRu*|���#�[e��	�iMb�3>��~H`�is��G6J��8x��N�&�b��/�6.�S 9�k6H�a~=3��ר�5�_ῢ8&�
�o`s�Р[���
=σ�Dw�C�`��1,�;����=�>m׵�2.*)/H*r@=[���&L*f6�ǻzZ��4�^��A��efu�{xR �f�W 5������4W8�7��.�u��H����ym2�1��ؙ�T?1�C$�`7X?��@�}Uq!L��8hV���-'N�h�ij�l��J����ࣞ|㩀]��5J����mGP�p%��]�G�l���K����iz�W'<�Y51�1
?�8�O�g�{+��<o0Fc�T�7�H�@돮�x)�]O��e'B�uvK=�*{�s�w�(8�P��l� �t��i %�fف��?f��ӣw��~��Hp�$�c�l�`�o��vHe��Ɯ�G�`"��B���{�F�z�w㿤�_V	��Fe����+�;�#�ςg��݁O҆�<�f�����da�`r%U��.�牊���0���.��U��GSEՑ��� \T���r;��R�PŖ�
?�k\�ֶG���S �� ������Zɨ/4L�m���{������&O�k ��W���(��-2B�ʪzҨ���zn�Xe�D5]�a0"�.p, �U
�R��Z�������Rs]� �6n)�L�8Gj^(�?�o�'����5F�y0����ވl(� ڎ_����z�N�PyŚ�W��.�u��!Пvn�L$���AvY����$�Ǣԭ�d'�!�e�Y}�1&}K��E;��c�Ó���V���y��-�!�����a�uN[�=���wǤ�,Xe-OtE��ɖ8B[r��[��4��'�~�*t�cu�����x��j;�����C�-�:�G�X��癭��K�-��o�<�YnS�.q±/����I)v��T6b/7�*:!d�T�!�������G�	Tt�[futlւB6�n3�U	�𸘇U�H�R�FZ��3��n����/�:t$�A�i�$ߥ������}B[\z�jv>��qц)�y�����/�׆} ��M].1���/(ɹ`d����2�9f��r��U�󆹀"�M{~q!`XEH��-W�(�N�a�59qn]��x�˙�k1��G9�VO��/�=O(bVV��k*Z�p���^.b��!+��cs��|�̈xW=�/����k���Q��K�T����d!�Cc���b�33zid�����C�k�Э>*���,SY����L�g�_L	��磤�^�o���+�B}�F�Rg� 7�X2V��"ε~6.�(��Z��rU���.�VD�O�o/���C���S�n讼�D=aނ�����%\w�KP-gɜ�t��e�������d�ςr���0�T8D��ޡ�S��b���'�c.k �?�B:�Gc�(�G)c�ǂ90��s�t��x��k�}Y�����Υe�?�ƝB()RW����tJ��wz�v�n�W��������8��e���`^�wӺ�F���g���T)�<�*��/vnz��s�Eڒ����-X�y�1�g��{�����U,Sʾ�	!��h����N>��q�|D��w�[���ɒ�l��pb�����W�۲��'~3����[?8��e&�e�J�IS%�Ko�]uX?-���Wf�ܽ�V'q���z�Tҕ;7���**���$�A�I̚ic� ��i����i"���d�j͔�_˝8RR
~�=�S����摾'��P�N��1���s�����Vy�f)�������jd(9�|�#X ���<0�~���lFO�L�N^3��ʆ@#w��J]�����T��N��X�Y4g�=����ru�J���>
.}�G%�����  Iгƚpo�HW�@�U�Z �4�s��o�u-0 ��bA��A��(Sd�(�v����]��3{D�t9I(���+�B��ܗԖv1�G<>�_����߳[]_�XX3V���ǣ���P�h�@���ɖ�y����,;�����㉋�e}O14"�i}���l��ç�:i�tm��Q������R���*�&�g�?������p2%D�iIe�J������)�DХ<��׭���h�ŗ��^�D�y�.M�>��2�mFB�ؘ�����V�\�P�me\*ӯeK�l�� ց>���l���%0�A̴]�E��!�A�ǩ��q��ҔU��e�b�#ZԸ�n����V�ay�l|.�{\x$�%�8���� Ju!�Z�#�"��5ج㑌��Q�����g����º\$����W�̨���$!�j��U���T�9�';���zV�Vnc�8S�q݉�ZG�t�K�K(|�ڊq������p��t?e�v��8��@JRT-��S��-�^��cPӠ�x��9�O��US1���=������E3<x���Zfqk��i�3JQ:\�-�7�f>�M{��ņ)�j�$�بČ�E�hɻ�u$\ A�﷎r�cr����h���N!3m����ҽV5�7�cNXDO��2t�r��ABd�B7�!{F��j ��#��D�:n�1����|R�\\۪̗e3��!$���t!4�����\m�� q��g"3��բ�E �V;	{���ItŃ����X����7O�3�-������0�����*_^�ꮊq5t�{�(��������'/b���pxK�vZ�*��[�����a�.����\cz7ͱ"�pŃ��@����ZXg���U��R:��ʉ�Z��&/HM5��� ��-���LX�Fp��~����7@�	���O�4Pm�Ǣfy��#�.\��}4�Ho6e��b�Wq>��kLlm5Ha1��s4O҄ʓx�0p�1�Լ6�В`��!�����ٺ�:S���3~�$^��U��֖$ Պ�)�R��DX���8��˯"L1aS�K��t/?��T�T�z�O�Ԓ_: ����	��8GU�C���-H�ZB���L���R��ֆ��NM1T)�Z��RPA6��]��a?������-�L���`l�痳@������w܆�]Kn�V�8���
.M�h�:�����%ڔ�[� l�:�������c|Y8���`k�K��w�$i��y_��&S��吊�T�t�&HHh��l���Ӝ��bԕ�4`�~@���6p�	3�!&�#�����1�$�������*�hFQØ�p��*�M�X�;|��0<���sq�Od��f�ɿ�A���1W�4}�^����J�!]�u-��7DN�V�����h�=����@?$�61�T!	>�sfp�6P������f�+�LY&b�]�i�@?�?���`��i�f��̆�!�ϩbS��]�~�̴"�_� �Z�6,��?��1¢�:<�aDw-��Ho̛%�u��8��f8Q�B���T Q��A1I�[�Tտ����ۏP-�}oyp!n�qb;٥�vk�M��*���-Q2��v�q�����ǫ��������<�6�,�\ґc!�TY���;O�\!K�\��gw��&,���	�s���d����hp�tC�t�]߀˨8Fy)��n��Q~� v�P��ܧ�p��rs3	�L�n
-+�l��k���
=���Gٔ�ߡ`�1���e�sZn5av�o�8��#��8��G�]��4+iPn������S�]B{�,{s�	��j�UڶL�+v0-�J���koLRo�i�0{;�Q.(���k���ٿP�҄��Oh�i���%h*ۂ�5����{y�6�9Zq���������:�{(�)ۛ�%����ᅡ�mm�9@�J�@2����3���
�O{h�蒭7�ce~<� ��-����ѐ �`.'��w8Ms+�~C��F@���U�0�#u��_��Һ�Uo��E�O>CXe�^������'�T'��e�^/C�.Â)Z��o�(���_�='V�b1�r�i�4w���̀���hW�ShBP;3���Y�=A�(���{��(�Yxg�|��P�Pͮa��<��̿�NZ�9R��L��	r�TǞ(�� V�?�~?։�Z���h����;���8^%ct.��r�l��Ili������LX�f8�i��RI�g6���{��
�5�b�����@���jG�o�.G8C��S%W x���D'�6�f�Q����?�� ��>��������T�L���h�U���=X������z{V@�8��a�����Fo��9�ƒ�>D?Q��H���S�EQ�CuM˿���M=�8��!`��VW��mV|��\�9�:W;�-���cW���*�c��d�B�����7ꇴ9����eaP��� ��.����
+9�P#'�~%l�|YD��@;���+<9}��w���X���g�>�����tB}�(�s��v��%�4���M���D����5>����_v^['`��2U����{��%�P����&�T�����n2@�h��M�s�|!��H�wb��z�3�o9�n��ok��]M����}����{e��oۜ���~4� !�J=�"�f&��P���Lѩ��E�t]:�
}s�9�&����������\Axh���k��/<�5$>�0ZÛ- `1�����^U�1����u�FQ!�^ۂ�x#�]��$dr������&��ȧ,A
׶�f����8:��@r5ʸ��9��k�r@�}��+H������lԎ��]A�U���GCP�EV>���Fw�����+� �'��z�n�^���֌n�5 �1lc5~�ܿr�,�`�Ҡ2�Wdz�$W歹�Ͼ�XE&�U��қ�0�xE^rO���ƅ$"L$��s�l�
��^�$B/R�Q1���?g��p����I(�Y��б~��K@d{�G����p���8e���j����ڂ �Q�V4M�x���|�MW=���,��l&8�E>�MB_�_\��I0��Swl͵2�&M<�H���'2E�U�s�mZ?�٨m5lw��A��X8��L���m�TN���Ȯ�כ��~YمnC�(�&���������Y����Nc�֟�}BS|���tdZ���(� �G;�ᄿ�_%�{�=��Iq7����-��ö�/����e���C��Z�A���_?
ƪ�H�"o�U���1��}�-z��Sv%�V�c�� n,B�#�J+=��S�լ�����voD�	&$X����:ľLc�8��Zl�"C�e��c�/�0�^YIZ%�dr�B�Mܜg�7�I;X�8݊�[����C�~�0띜Ԅ�Q�kS 1�f%�,���+M w���g�#*��q��O���B�IfИ�&b���rv�t	���C�i�xͧ��g ��l�3��T�0������t�0�l'K��,4��K�d���ՏJ��ȧ�5l.��c_P�T���(ņ���F�D:vԭm(3�����D.�5�vpE��m4p���
=�v���'�4u�� Ӽx��""@i-C�q�Y����jey�?�2>[(N�V],n�<��3��
j`�?P�}�h���A��Ħ~���{�M%�l�#9A�7ԅ��y���[	�i��u����v�4���*N��6����_ǫCb,�<���2�b��/��&͖������Wq�z�0w�3�'@��jwu(>C뀽���Ί^�Ԋ;{����𷢊��r�z��/��;c�)�:�N�\�끡�hU����E..��!��~��A7 L3�|��U�R{G�d���,����u�����~�$�*^�4�wGQ��^@��ދ���*Pn�� �����qsp�	es�!��ҡo���>�xc,b5� l�7������ÖS�b��Z��?��e���X?��@}֜W��r/	౱��ͤp,� _5�̍����!s-��3������_[�H��SɃ�1�@� ��GlEF+ZA�B�P8�D��-�b���#�������gw�2)n2T}�Q�{֠b�"�mDl�zo����K��sP�AϜ��W���e���-�aAٻ�;k-�6���ؒm�1��؏������?]�O%n���tDS�K�?�+-���3_ q�a
�=U��@��8�ڱ�dŬ*@��#���@�s.�F1e�>4���i�<�ŽBB�)�5�Q�)��%jC�A'멅���]�������M���rƙa���
K������+��G8��������m�v�Đ�%�!��'�du�Y9���,�m�Kj���q+�|,@����7���.v�3�*�i�1�\�p��3ܚ�֭��F
���)[u#�訬W���49f���"3�.�6.��G�`���8��-�j2��1�"�ȭ0����59O�%1���G ��yw��M���=�1�|%Q�(y^hօ�e!	/'Ơr#}4���> ����R���w������UH�G� �$Ng����p��{���fԊ���׶�������=����H����p7��	EN3;�6�Jd<0�}�Bu����<�H}�� �C�YK�l�> �Z�3�7���f��8�]���`i�\.�P}���>�I�S�k��B3.s���� ��^�5��6����o')
�ѓ�e�=P���{���<Ӝ�w��NN�9m�����vp�m�m�v����]|��`Tjg/l�%!��^��&c՘/377Ȅ�!p,�Y{d��N�T�M:
�`g�oc���9h6,zˤ$����6�C�W���a<�4A��@��c$K+k�2���y�=��p��L��xƿQT���7��G���5�d�7��8������)xBܪ���p��-W1�]8���4��S��hW���
{��K��h�����&�a�4+��EB�S�-|J����]QfU��r�����/��x	V�D2�I o�h�y�6�Ѹ�!\ڇ��Uc!W�'�o�|�^W�uu��[s݉��j\*��{B,����2@&X�+f¨/���A4����{�Rr���ģ��	�H���ט�AO��Օ��Z��ZY>���#�F��H��k�(C�C�x-�@N��%��$���oeX�������5:*A���R�U:�X'{����ϡ�}g�J�cB�	c�$��##�/Z�9_�&đp��h~a�zh�r���z�j�v���x"����|���Csa�P`��ݼudfa�Ck�:ڈ�yK���,�Sx��Φ��@���z�������7�������Fb.���p�=�i��3ĪV�P�c��Հ�Ot���*&��B�,�4E��^��I'�ګw�Q^0H>ޔ\�*;�^��>]�o��)��A|����C���� <�`M�[e�Tqچ�g�����&-����3=_#
K���Jz2���K��&�G��̍�1V�}w��V�e�{��K����]�]���]�{a�b�?�g�%�6�l�ͼ�\�������#G���JU��r���A�2�;�~�>-H�Yt��|5#�/�+�&i}shŌ�mA�x��`�7eE��ǫhKn��C�� 6�@�yc�_�8]^��'m�g�da4\M�_PD̑Y��_�~�g(dv~��Qf��_AO \��&fb�\�e�mh��#I;�ޭlR�Q�����
�Lun*� >��b�"^�D	�����f&�N Մ��@�sЛ'�y��FY6%N{zs�).X���)�C6.IxM�)e�?������(��n�������P^ayV��$	�%��O���� ��y�N:���J���³T -�r�C\�P�v��.a1�*�#��j����_�X�4��D8��o��SChß�������C��!&�@"�29���f�T6V��S[��	��e�����	���[���y:Ҳ6����ˣ �$|��c�Ή|��T���ǃR�Hb�^k��[)�gd��ļe��Q�Xf@�n����wH0��T���^X���&��iM�#��>s��P�-��x#eҺa1J*�5E;����i9�'�*`�j�%��$MGZ�n�Oa?��g��;�G�z��Y�h�$j	�7e�> ��򧭀��}��Z��rp!�<�~�Uzj�
�ȅ�o��X�J��,<\�#��b��E$�d���Y��}����^��Ғ/�a�q�� &.z����#�.Ŵ��������M;�_�5��ĭ�gR�m��6��c�y4��N0��ג��E	��)Q�r��H�������� �y � tKbk����$F���#ޞ}<S��_���ɭQ`��vm�����1�$���C ���5�Vu�1M��bA6uFZ�@[x#����d)�{"����]��]�hh3���y�����vAA�Z�=�ȶY4цHN`�ՠɵoki�\�V����8��O<s�Q��C�7ܰ�t���(~��N�̰�ލ�T�'��7A^;���+��O%'�"L���zv(h<����~���1WZ�̛�5���w�%:aa�ڂP�m?�~t(/	1���ơ���r�ey�д[[@�\�T�{�v�:��{��Z�����l��	ِ�����KiFE%PmS���碦.�2�H�s�j���z��o���Ih���o\QqO��rAV�e����X"M���q��:���&b��R]�GDu"K��0�����6�c��@X��XW2]�a��!ϰ���Y�s�dZ�;�(Ӕ��M�Ž'���0e�7C�7$�����!��c>q���d'+=gG%��	_����� ���Q��U,,2���Aڙe��Z�T$��_l~�^�$Ӂ�ڦw���*1��R���?�9�{��������C�����h��ڶ���pꊓ��*��Qh���2ҫ���Z���,q���*q
�,�TU�x��
�%4�gnB�E|꧀����:R�߻fa�MЏg�*8K�ܿ{�:2Izvx��ȥ�M�#ۀ?1�b��eYv�ŀ��1*XSw(�����4�p���e=���@!�%>:���#y�����Rq��@}I� �Ƕ\lA���Y�M����, �~�D�H%��O��m�YlDw���]&{�b��q����!ܘW�C���z�3�z���
�/;6��s��RXƪ��;(����Yc����tuo���s�s�8r��6ci<>�U:�ǳ���:�C��Õf���İ�_m����8��}�#���lb#����	��a�C���H/��Hj���[�Kל�"��#<�_J'�΀�D[/���uߦT	#mvK.X�;������3����;;�e� �;�b*�~�[_km�gvT��E�@7������h� a͋^�7�7�>��1��� � �����Zf��)9Z
�>F$����/7`ݼ���^yx-i���5cptl'�"�\�>ֹ�m5��y�ܐ�X5,�������ڵI����1�+ܵ1M��9b�\�`$�������1�$ţ-�����5�vu��8�u���i��%�	����V�3����q�Z4�� E)Hx���^���D;��W�-�q�'����L���[���(h��_�*S,[S��L{O��m; :���Pu�T6[���q��O<���L+Cu�wR�S*����(H�8��c�r�MPS�F(?���qJ..Y��G�xI�ቨAiXrP��oۂ� �����׶�չn���HD�*#,���o�\�����PS��:%p#U�*2�1����Y,Wu�9�haO!�l�X;�Eo8����P����3b�R�q��z:����D#c���blI�w�[�� ���x�̓îŊr��u"iqu.�e�ٷ�9O���1Ph��i2qwL��[ٌ1ĸ������������bظ�[��΀�˳F�2�eG��-���t;�VVв�&�ۊ{�E0Qg)ٹE�%������Y�1=JArlZ&V�e����o�	7��m:��]S?&�LۉE�N��������d���*��3��\���NĂ@h
\�栌��@D�~�X�����B?�w���x��m�o��x��3&�b���3����랁0�F��AY���k���P�8~!�R������N��5 �X7���S2�J�&1���C��?��K��ow�u[+�a�8�xA4�ٶ{��ژ�P��$ESG�	����n���X���7҉Iĉ �m�"H4�:�@x+��`;|2�e�%��eØ	+��F����m��^���|h:!Oh(�4#��"-�pH�W�*?�oR�����R�y}�z�0���~�1 #��� ��J nI14	��sj.g�>]Hr�Z��Ǿ�0d>� /<�r��/�kE!�ox� ?:�X푐�b�~}U|�,d��d�5;շ>3�X�n}�����8��e�p�X�1m9>Ŀ�1D� ��Es9�Ц��cJ��ў6)>�Cϕ]���;�%5���� (�gJlY��2�
�ӄ��)!�@��B���C��D�IGZ��GC��ܢc=�su�.(j���l����PYҽd{�w�PS�9��9r��ԃ������㴻0t�m0/���F�'�CV�A\ x�{d�9�wn�!�.1�?\��6��3�;1_���Yj���*�ql�՜e������on���{T������<w��~��r�H�ŧ%�+C��Uu���#�c��pbC5��ʵ�躑i������e�՜�|E�))�+L��
�R;���h7�>��ȓ&V�aϑ�J4vϼ�������4���̟7����Q�>g%����N"`% ������!�v��om����br��6�p�-y"�f��FO�b��h{��n�A+�,Z����y��4��}�y[�yl{��(3ҍ%C�ߒ�v�#2g�ږ��<� "Gz�n,a��շYW��H��V�5��޳DԔF;n��y�܏<68�SJ^~�
$�sЉ��0Rtt�E���t�\ځ
A�5���K�0S&P����� 3�{���@fv�U1�؉�y4�Ahw��s�Z�}�T�bj<c>�P�G3"٥��$���e��Hh>�؁^�i��uL�xg88h���'�/�԰{�������9��+�5~�_��_������]t7�6��7�A4�"��#�W$+<#�Ǫ��^`_�J���˼s���v�?��\�HK���-��ܩ[1CDJ�;(o��J���!'�Y�Qa�4��/ T2K�fc�U����H��7Zۿ���Q�'���σs>�~�-��2���R��>9F������{�1�iLsT-o_�������EkiT�^ �/�Xv1�>h����Z���]S��o2��}.�U���9��G�Č}嶚I�\�j�Z�<"-6j����C^��`S�ة����� x>w^Ja?S_3<��o�}�r�QH�0��!�{& a�>W:F�e+R�xN�%?e�ʳmo�7g�	?5���y�Ĺol�b�����M�F��)Hf��4��V+�=��v^��^==ߞM���Q��Jb��e�g�h;t3VO ��Y}K:������NU��Z̒�v�k�
�� �5���9���γ�c��ϛ�Q�s�-Sh��E����������+Rc>[=�k�{ކ�@0�0��{)<cv����Ո
����oR�jGξ1r*]*����H��8Jz����D1��j��^�Ʉ;���=)#�u��0f��!�	C�˸�N��б����7�i��;���u���uի�A�ݑR*M7�χ���uZ�,.+�
��=&��#��?�\k��?���`� �_?Ϙ2�)0R��.�QQ@�Uw�s3�l�fϻ��Qb�����l����Q�esԖ�/��P�k�����n�]ڋs0`�7+(yKK�}k-���U��򤖒���<���V�Bln7���'�hO���(��@�$��$�����P�
h�]|��2d*[~ע$=M���V$�O��R$�d��&��Xx����Cm;�~1��������+�F�Q�OL@�S�E�
�Ӱ��!�|�Wl��.�N�=�SǅIXw �^�b�%�8����2i���������>�=��?��N����[
g�p��_ �*�W,<��xw��A�N0�����S6������(p%�v�C#.!|-��"�\�sm�xA�%|F�^���Y[�\�v���'�\��eE��5�����J]D�d�*�R�gu��d����>�l HG��"0� ��i!]s� J��f��΋v�౐!*&ɶ~��&v���h�G�Ԥ<��/쬐9i�R�9��b]���j�ĕ9�"�yhD���R��]��{-��x_��ԁ����L6���!�A{g���2���/g�2�@�{ny����Y���\�N��Ƶj�P�� ������m���ו��H��>����N�;"��m�U��2�Ld��	�Mti�)�u����R��H§
��x���@���O˪�&Z���-!{��#1��.K�q�e�b�,� \��;� �����u�5�����,��'Ǔ0?�׬�X�I�D�>�M.)bw	��S�������-P��j$�b���3��z:#!=��d �̗|�l����,[��byIT�j#~���sI�$݆��)�]
x�J��ק(���oж߰�ƫ$��F�a��S�L�)<)~�w20�ӽ���b���"2#(OZ���'v�w��o��Z��ġQ�6 ���[��#n1ݨ.}a�x��g7_t���?����r���
y�S~tH�!���ֶ��l)��g��������.�B1f��X�{�~4T�p�2ۏ�}�e�"koY�d��x^��u��쏥��ޤcIG������~�I�d#�Y�6��]�,2�9���/Q	���%D!�7��z�ެ�b�����n�>��o�d��$�U9��#>���o���dw2X5�U��C��"�KA2�U }���%N�b��Dz����@t�U{�oo�HF�?��aȤ�6���瀈�h㪩?��2C����H��2��~��\�Up{)F�}����V�4���Є�ͮ�Q5�q z�Ad����S�]�
蓌�"��[�V��qʛ�Zp$}-�ƞ�t�G�Ka�!\DR;���2��O����@�2z�b��y�z��]dcU����!MaEW�?f���4Iч�͠^&W��t`�|$3�$�э����,�C��g�_*��
R�.�I	���PN�+i*�q[u+M�K�c�z�+����7όN�nD��m'5���H1ޙc�Xl���R{����b��_M4����E���?/���+$��
�7N.�gƗ������^�ʿuJ��E�s�����O����yM�NK�����i��-iLT�:%�������I>��<f�:�Z��i󌮖Ct{����cS<�?:5Ut�p����\7�����a�p�U�QI�|����q��a���n�%Lj�ϋb�S��'M��߬���	mN�w(���'���sF��T��f� �k�ܛۚ']��DӸ(�
m���4�ݞ��Ճ��E�ok.���k8�Ŭ�+�!W5V���m0�����j�Fj~�,�ʴ$�֬�|�mJ�����/�p��нm0m+M\w�TEHuۡ��/Ϫ����`����q��R,�/�)k�Z)�\y�$�hV^N��Ԯ C�K=��юl[��q/��K�Qlzw�@j(��2)�K6�?-w����f"]�Q���5�n*�( |����r�Y�+��K)�6.�sVhО�%��W��%���T�O/��+����:g9�O_���~�`���oG)�ݓ�J����*�b2'�<�O��'���j�M��*"��39�y��O53��ȃ�)�pЪ��{/�o�)'��n�gZ�k���$1�Cxr�qp�W��P�6�X�����.
ejJ����@z{���������$9T�Q�X��#��9�t��ά���R�|,�;(yu�K�[^�*�4�F��mʐ?.7�|2�x�N��Շ�(o�himBǔ�D�ޜd�uA����V�-��*d�����_���p���7��D<�.*v8� ��4. ����v��^��VD�k��,Bb��pJ{��L��@]�q��	kH���&L�@~I���)�M��Ԑ
k`��+,�//��R�nŠ���JY�`�ŷq��t�O��ސ�C�xn����p����?�ն����kE�H�$
���K<at����(B���M �BhUl~	��&����吧Bٛ7��.<��2�:p�%]=�D��7`}�:gkJlL�m ���/�p�qQ���}����������i��H�i�� ���W`�����;�
�z���d�=���K�;���Tr����Xa]N[�O;���	���'�1�5#S�U����i�(.{�-���a�gM�s��j���m=-��8�փ�f=��((�Gb#��^��9��]����!P��`����`��)��ZsZ�&�����Wr�A�.��#:��@]L�N5�ܹ�N*r�iQXc��<�UiOH��o8C��4\�$�����x��0h��}�S��Vk7���)_Qq	�ٜ�a}F�O�M��
QQ���E�YK�08�
���ˉ=[�N�o��P�_�K�ρvr�/��o���>��O��X�x�?��i8(й��/�x��mj��/��zeu��>�sK��%�z
� 8���`�<����Ze_#�*�.(?�|�e��2q�+��aV3��1���a
n�٭��lA`ێ����$�C6t��׎�l��}7��Q�.���E�!�C+屵mV������w���@]�U{�>i�WC
�5�x�<�,���ə屢p��)a&��}5O�!W��L��Q-oo-�X�� �,�\�01uuvl�x��+l�N$c[�I���*���̔�xQw���3�� yi���R�\~�������p�u�V'Po��G���B����:
�gSو�r���+^t�Vfm"�y���E�c wq��&�}Aݻ���tz҄�t����jY�[�`H�O�m7*`�Z��':� �x��0K�Ż�#�E�O���j��[��G��� �)ք;�<����m�vD�Zg�'����q�H�4s>=�G9��2�4�v�J���\p�N�a��z$���2��^�W��G*��6��Ok8bt��q�F�c34��� �>ue��C�tM��e���*N�Qd�i�!Ep�u��v�f-ŠrF�r�)Z��d�)
��WA�skZ�=2���7���J�'NO���<��?'�`�vHu�1������'�Aْ��[~�5�^�Y�e����r|L��j\�s"�����`l!���v������)go��,CR��L�Q/��rsE�c���=f�[㓢��􆹕=�]�DF�=d�҆�K���B��qZ^f��C���%���i3ܝK(� ��18�
���Ej��<cN�K�ZnU�)��f2.<���h�fb��	=y��,�KC��9��;�G���s��r�8ҫ�E��n)/cvN�Řϒ�,��=�,)
α�A�T�8N���Xp�\�.J7ȹ�  1�C�u��%#uH;��$� xJr��[Q㲓�o��7�y���PC/W?��)!�i�����&��ʮ1S�Q��?vxo�w1�P̧*�a�~��=����C�ޓ��}GX��􋸾����g�v��iP+�AQ���s�5H��q}�4���+q�D�?�D+������ٔ�F���?4�