��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b��%[��$~��=�&��5J��$��_}l���3���ed[ꢂ�Wh!ڭp�>{me��Q ${F�e]��x+|mj_^Θ$�	�� �5� � ��1c(�,�t��S���8Y�nޛS�c?DkCK�Y?ʖ�D�KL�$�w����>��z�`��Rk:1��/�bZG�۳YzY"nD�ʩS,*톈�_�� ���mݻ��0LE<4RD"YpAB�`V7����o�1�4"_b*�k�Bq5-�/� mʙ	0}�"�O���=�
#��!�j���_Wt5 ���z��.�P(zSH��;͇�n��K��5��e�@Ct"qa-Y_��]���(O&���5���x~��m;wZK�g4��{���tZ���4�m�,�k@K�������0�u(��8��ec�nI�������R>($�����&��Z��B�%*�)O�|��P�l��/�����Y@?�U����j��X�x�dYGD��L9�zb7�I���J�+QL��ܚ�K�e���S.؁�*�w�v~�_P�_�(�D�Y\=�>;��7�g��S�~���̫�/�4Q��ݯ��a�E��T�~��gY��p��0�4�3��>zC����6
t���n�0m��g�
$QV,�H�'^;ה��ʲ���<��U�Z�A��/�N԰-����?LPr�r.�z����\UoWTnl���R:�1{8�K��jH����F�V��6�ʠ��*��Ճ�ԕp|�ܙ�4�m� nm>q�,*x��O����]�����o o.�˗ZƄ tZ��Re	&����CEh����UE+���Kv��%��f���ˎԲ�-���bD0�ޜ��L��F�5G/lC�p��K_j����Q��O/g�T́��0�Z*�ix���B~�x4�􆔗�T����;*�,�G�����էE��.�)�%��sK��~�En�a%������qU�o��s�/:��}?���oC�Q莰
Š7V92��E~��K��P�vĚ��*�K�'b��]G�gh�'��H�ƞ\�P��I:�qDҐ9u��`�c��D�G����#a�����C���zQ��Eq�p��Y�J'�[52"�,XȖx`�1\�B���Rt�O$G�Y���2�,��ڗ7��VG�5L�^x�>��>�k��3�[^������ɘُ}uz�GǴ�ʷ�?�y������Cf;|���<a?+�6Z���B2�-�pD�6,�.	b�������k�ݙ������x����KM���`gR�c�)8��~Uv��0���l(����x�'�Nıϵ$`��7�q&�ׯC��|3蕠��c��a]�*yAy����){�z F���Ez �Q�P,��;U�4`}ԑ��e}��Y��W
���Zلr�D���n3����{bӡ'9D���P�����6=mF{�灃z���sR�t�gm�X,�X��|o����ӛy1��ׇU�UD�|�j:q}���*Px��ͩ���hV�Tkj�J���;V��>����
:��☠�$��ɫo^Z�EM��iڈ�&7yQ�Ə&����n,��R�� ���{�BJf���<��{<0E�Z���Q���b�L�(�;H��2c	\R)s��U��L<2O��8?@����G �m=[��D*۳׷�̾�"tu�~g����:�0X�e�
:����mg�Tz���?_�G�v���z9�~/���FF����0=z;�
\�ޢ����J��m�֫H|2�����H0̀y1?�@j{�Щ{��;Dr�3΂�cnO�����hφÙ�VR4�EG�PJN���rA��h"*R3��|��۶6�6��W�LZa^�I�f�2.N+�y�[⣘�Z���=�����cp"b��JPZ��w._��p��T�g���������;�O|`/�lHINZHA��j�u��0 � Dk#]��?�.�u��d0����H�����X5`YL��j�C�p�쫪$Cq��.��!��~w�I�V�����X�fQ#\�}3A��k!��A�6U���|Z9�'�_6�~�d�'/�=p���9i���c���NT$���3�8��8z��N��u�K��$�0��!#�A�	�����O��ͨ�ԒF�����f�M�4dM=u�רۭ���6�8qƲd�����a�l�Z���t���69��os��v��c�h�H �ۚ6��c�vэ8�"������g�8 jw���0���Wq!/��M���HW.�!)Mb{'J�O��Db,��Lh����V��`�ܕV����B@�tT~�s��6ha����1:�tf�5����6�.A�|���o]�>bb5���K��z._�E��'� �\v�bV~�t�F"�!f�|�� ��I2*�m�����C��x��,�I��Gɇ�D|%Hb���Nդh�1b�.�OC���0�Eݿ�2nћNk~��'?Ü�	���!������P�J�종����
mx6[�eK�1�����&�.�b�HQ�v�M��2���[k�?�t^^�(��.:{��~�k��=Y �o�2����nS$���W�]߃��;\	J
���ֺ��͋n;�M3�R�L�S��q�,��]�%u�Ozyem���.Z��p��$uEu�ǀ2��dt��(D�9.[co�ʾZ��V ����ė����;�m���=�>��}���&O��N�AT�ڜR�uS�w�(�����B���S ݣ��>޺T��6 �"иD.��6�ts;C^�m�-M�l �˿��4�r"qj2�">+��Y57��x.�!���w0��m���BsV�3Ȁ�ucf� `npn�ԘI���ft��gG7�_�J>�x;�g���t`����T�E���N�p��z[H�
J�����c��3B��uK���0�,�%�I����#�;{]'�_��ȅl������*W.�,��a���V��έ�t�X�4�xT?&�A�Ë0��G�<Y�Z��r�d�L))���@�&Y�Ð!J�E�t��^��eӜ�1T'���c�Df{��}AΎ_�2���O�	�OoT���y���	�w���[Ä�P`_�E����RleC�n���Fa9�y�i&4���ܒ�"�����=��rzM�����:����N��y=0WI�K�����I�8ƾk){Z�C�gE�ǭ�������lHה��	��*��7e}��E�r4�.;��b��Ůx��!
�'p��c�{�����h�����^��a
�2��T��r3��^UN��ֽ巔P�/�>_/���Oc-ĝ+҆�����~�UC���|ϦoL��aS;s8��\&P���\����3f��́�	wo���MùNE��k�<ңI_� ؾ��>Gn=+ү^XĚ�<�S�i�����@��_A�-�3G2-�n�=�,=��NҠ������$3{W�.	�Z7���ŬUQH�^M��bo�.�I�K;��8ŽiM[�u�[|�`�p%p$���R�Vs�� x��PW�j<'h�?���懯�����Z2a�E�����n���݆��᪍6>a��K�I(����T�!���!�e��^+���cK�p�3P��Y��}م��`U:��<@��=�T4B�䀉@��
��z�Dd�*���ԟL��Gm�^��}��%���7���n���_�n?�eX���F���a!�$�Z�Ú�R;bp�>��@�3���D
�R�l��[� t7wå����K]��3m�sll�:���g0�%��d���d|4a���ƍE�-�;�D�@�u��ա �]n����5��u���J��ꓱ���/���u��f@���@��_�x�n1U�"�R��כ��!�5�$~>yږ}r��[� �@[�1�_��������
p�:) �4�׉n�?�:�F�)
�Q�f�Gu���3����}�U�����]��7�:�؍Ot�NGp����M�w^!�_��@ɪE������w�s��mT]��裸�G/�~�t�B���X�L��}�ï]:r���.b* ��L9C���󸡋���CU����D>��O�k6A"������o;�KɆR��P�H���aP?1BBq7`$�/��9���7�n¥�f�H�8�\���ƨ���
��C�ksF*\����Is{�q*���֌����+A��mO2��|)NA��p�^̹T���8T`�!␕Y+�
�"㍸�
8�Qj�H��D�7���\p��aD���N�ߤ[k�].�Pa��DN�	I���jѬ��޻�C*J���ܲl��VɒT0���4��0Qn}���	}�f��m^v��-�����*�zKE��ٮ7���G@V{�iC�ͱ�6v����eݲ>S�~�vwj
������F�)�YEÖ'�B��3��0��6�E�)��r���L�0��]F���xr�5������v,ƒ�4!,x������\�, ��}�!.lB쾿��V̍<�e %�!�tuny�D�7i#J}+e{5�g����u���3�~@�����rs�5	[)�m��v]��W�m;-��X�~�bPƸW!�O��kKS`T�t��#h�D��e����z���hUȽb/�ک�Vѳq���H������ߦu�rG
�fKDz�o�{�\����9��8��b���e<y���Iz/��G���w��L�C��"K�/�n�{�w���殇AqT����J&P�e�(�%�O�T��q#�O�͡���4���e��^~bF9�]��H�P��B���a��U���\�XTp��nNҪw�٥z Ð�,גG�"�p
�,.�����p���0z����X�2�v��㦥��D�`�'Ct�@ �,)��[5����r�T�>Cx�]�#��g	"M	sxC�!+�f�y'>�g��w�#+�g5��)\K�{3����|�w+�gSA��:d�@9�s2�$�Ե���`_Ղg(�,��ĵ��ð;'l+��.���or�АN���h�G�nӡj��1�P�V�f��z�S�(���@��M���&����gW��*a�H�!LX�}�5Gn��kd9n#j��e*05�Ĝu�1�F�N�Q��g4��:d;���X~�^�k��Y�"�����JJ}��+�&P�k;ҡuǳ��VB�ɃR�ا�4T٣a
AE����"5�����I���5�`��l��7iEW$� Nkt���݄Ձ8!2��/����?̚�i���y�i붭T-j����fP�Ө����e/����`�]�}ƍ�P04.��\�k�ӝo��� �����װƔ���T�h�:�]! 枡���8m��Y��P��͢i�s=SLW8!��GZ����&Lg8���V�x��G}8H��٬i�M������<_���]�-���a���݁��9�&�f���y��H�*�hWk���g��!��y,�d��"�ȕ�bi/�D?�t�8�W;�aG���F����tq�v>u"BS$%ΰ��PS�6�f���0���]�Zچ�R	X9 ֩ v����;R����>�2�x��dݱ޴qn�yv�B��+�ze���:���|Q	�/���	�Tj�ԁS.����Cn\��l�x-��-��* ��3Ş����mX�3�
"�3?t�hzڳ�|�o���2�~Υڇ���,2&��x��XWP]��@U�f��;7O����KT� �_��^.3؅a+�1@��'�����w�\i���^��ә��w��U�<����A�����cH>�Q�R##���s1����B���SNw �Q���1;Z�M&b:
7���F�^��Q\�}B�==|�眧}�ܡ�"��R������=u ,:�'Ý"���t��Ul�ֶ��-X�R�����c$�HtB�d�Ӌ*���rN~��hR ��	��@�خ��r� �!���f��+~ͭ�I��c�m��᫦`�1N��W���a�u�mC4Y�t^�/��ȩ_�u~�x$t�~�;һ�Q�o�hq-�Y��U��j�$�u��*�����<)�$$��4xa1I����z�oU����A�߁�;�=�M���FD�O(�������:A�/���C�v:#n��������_FȿW�j�x�V�v��}CZ�!�3ZG�L"��C]�>��N$K6�v�:2 Z(�� �PZ!(RJ����̠}�i')Z���g �D=0��J�?�^�G.Q4M��{��3���&�zI$��?�
 y�"��Z4$'�՗�N.)���R�p����"s嗆�"��$�
Tb�|�Ί��s�Gg��"�`Ț�ˁlL[�x�DUR�*�l�oj}�:u}ϻ����Kg+���7\��|1q�$���>����F�"��<�o�����٫uQP lQ��~�)��z$�y&�:K�;`OR���9Z��o��E���*�Q��{�e#��Z3\����OSlSvl��W��g�?�V�]"�74K�?��OP�tk$w�{��z�/{����$��例Ju��%�$��u}��Hs5�D��nH�H�Fj#����N�F!��P��x�,�8�o^�,�������/{�6P!�;8�z�Z�*qq<�E�P��A�%���`$u�͘{�?I��>d�c��J4c��S�k�ٓ:��I�O֖�%4i?KʮG(�C���e��6!�г�ﲘ~2�=�%�6�E�j�ܾ>��gݽz}���?4�S�Bux�;���~x�j���}����h�5أ�^��X�>~��x[PU�Y���M�#�^V��w9x�����P�V�W4����1���h�.0�е��+� ��o���j�a����̳���G���v�O.#J�xL��U� �8˱��m�C+���4^�� wv}�؟9�������W��=?���"����Jf_DIR�p8��yĘ�g�e?���t�9��,��'�
�Y$
s�j�0��ω���Q�h�8D4��[^0V	5���CE1�ӖMĘ��t��I����s�a�7��}m�+�0VƆ_���Kk��/B�& ����
g�P�ѻx�w�F�
���I���ܸ�q@eQJ���K� �3�w�̚a�x)ǳ�#��Ƿ����7������z�82C�EH�;�������6�jB��R^��p�����v̠���|=!��lvB+���<����ڷ�	i.4��������*.Oi6v���fD!Lv�	�OJg�h�j�y>�}��ښ��9�>�2�L;�Ec?62�n;ϱ���'�ɿi���y�'	1�W����A�v���=�������m!s��&q�rڰ��lA�������J���;��;�i�a�k�gf�����wJ:/~p���~��_���:��t[+� z���I�XD4Q�4)�a�fK��0�e��1���US$}��{p[B0��
��:;�Y��� 0��ʜ<U�.}Kw	�y�~K	cv@g�[��x��
�xf��W�Q@���g�5�z�̋��Z�gF�@\��^I.�|�el;)]b�Ɣ��Y<�<���۞E�@Kr�w#��.���EuH�Vٞ,T�̆�V����!+k�I�,��l߲&���B�W}�tk3T��4#�B��#	N�������M��I8`mT8/?�%���A�,��[�8�7��ԇ7~U����uo�����9MK�����gI���C�x;]�P*3D��1�It}��������Z��4f�͸L�n�y ��}�ٷx	��/�T�.�Yn��i? f���E�Es�L���)h���3�q���� %�r;2y����> 86�>��8��~��MJc�?h�S�a�<8E@t�r٬�t�I�����W�k�����E?Ė��Hg��zn��q��y%��4f����چ��ޱ��$fR�Z��n�g".���TSdj��ꀴ	ľ4HI�~�]?�p(�
��l?d$'��[X��B%� �DЈ�/�T�m�}�!��2���ά�
��YP��z�FX^���p׼`>���	<��:���:�(����I�3ps�-3�r�O7��fs�h{���ܽJ:`i��5��M�}����
c۽'��Ȃ�ژ�]�9%�MVS��饯C�ф���dr��EQ�ε�N
'���aUIrn`�r����_%����4�|.����9��{���,��nҕ	/���R�S�#�ms�%nQO��=d8?�-PR ԻKR�g�2����ze���2-=x.��x�g�8Y[���)���L�u���c6H��^�p���B�|��A�aG����w��}�I�ź�h.g��Fx+
����/�x��z�/����´
��>�^ZZ�?e�ry4�
A�
�#��f�dy��Ɣ���?�j��+4���d�.%%[}8�x^�8CTsA���X��J_� ��cf)K0t�R����8�|�.ft��Rg�#��8�?ǒN�!Z�-�@0��I�Ā�G��:�2\������.����@>&�ҽAU�; !��p����s��K`$j��=Q4n�k{�traW@�7ݩ�ߛ�΢�6�pA�?�c�����Q*�VH4�����9���JB�!{��aKj��T�����l��1���6v:x斺�y3k-\���y䚋�}s?=0�q�8�h�j���g�"�x�B���g�| �����d���@Ob+�}�G��H��R�4��~�&�	J�8��0�H��zN1GF�Lt�Aa
#��G�+�jPpm�ˡ��w2w�r�&Ч�=�%,��?�HyFC0���$j"�X�Ɵ�vߝ�>��9ݹ�/��ח��C>ƥEN�ˁ�7�OƑ���{��ܒ�e:��m��y=8��Le��@�c�ٰ5�ޱz&�(^	�*)Ha$Upx1eǉ�O�*��������S�R���%�RIj��v���|�F|&�.����k�W{	;X�����W�_p�x]|�ҵ�	j�r���ѬJȤ�FҽkG��䥎�P�y�оIE�1d݀��p��
x���ZL�Z��S(�e�Gu}��A���T���Ż�˧��c+��fǎ%H��;�3����xr��Z�e����WC4�M9A�A�a�E�P..L�iMI�a����H��(L�<�a߱�YY�fFl��cJ�5o����ֶlY�DbQԾ�~/��6�&������arvȌ/+��N.C��H�!(F��� �
��Cy���?���R�z=?<E��>���ގ1�<Pp�<�T �O3�*u����q�F$F���.�K�DK�����5�x�'B�&���jS��>�U��;���o=+���P�k���B��,xL�	9o�ߎ�T��$����.q���B�s�]3>��цX�У�Tu��yBw�m���LܬMW9�"��;(^Ƕ�\yK3/o�B�1g����/�N������a|��Q�,=0�''ď���|I"�W��D�o�_܃F�,~	�f51B,�yK ���G�H�?ʽ�ӹ5]w���Mݵ�d�`�;�0�b?��K��o��ل&��(�ڙ}0lԱ�ʈ�,��((:�* ~СP���C4�cQM3HߤO4�
���ѱ��˕�_^ZI?Ø�_����wQ�u{�n;!��Įg�V�)� }��lƛv5b�3ba	L<�R�{��W��i%�N�OIhw�V�]��kv����2o��� ��B�a���t��#�;���{s�m]H���rѪdz(�-��hG�YY�Ԕ�ʌ�d�t�{`L���ƌez���(���y�SX3�|��i��u!��W�H�-cm�+�9�-��A��_��K�f$җ��L`;��i�q��h�+���������˫��Al��!�����18���p`+-�2ƕ=���)���˯m�Yn�<_G�h�6��,XӘ��[I�?�|{���evLo'&�
P��2S��'�nl3p���j��{�!E �VL,��MDB�ՕQY�;[$]��u��F%�%���ܫ.7���H£�����i4�-jg��.MލvI� ��b�'��s���IIۈ����m��9I��}�+�j����7Ǟ���Xr磁U1u߫�؀�c�s|����8�\rd�K-��/���g��<�`,<)��*xy���׆�\��� h�iX*�P91�h@Qe|��ݘ0�}������P	��h��M�ύk:��Ym�"]H����<��X���[N��h��^�!#]0i������1m#fN'˰�H#�׃|2n-��bC�{K+)�\���(���n'������}C[�ږ������΂�:�_�I�;�9��f"�&�S�!�c�Z~�x[��CQp�����S�`0����B���=�3qDA)�nE�t��ʆ~-�5G)/�a�X7>NN5��Sڑ��+�S��+C;�BJV���ƣvy��s�$�~��|UaD�J�Ҭ���"k��3�����������<�G��O:�$°���g�u�T{��H?[��lo#R��9_J,Ë;�l ��F�a|�5J�"��2�N'j�Ï5�y���D�B���a}��ܯg�^>i�º��9굽:�W����OG��l�R�\b�0�Y��aG�y�O�^��΃e�p �(��O)�aT�����O���d^�$}u��4{�w�o���7�R4�+e]�6lLQ(���1(0�:Ɔh���[����:��� }P��NC	'�M�[^��cN5͊{)����l�g/���M\���M��j~�)�躣��9		h8�O(�l��Y��w��ԈsIÏ�0������&���̨��+ *Ra���D����.��_*��cH��K�;c(EwS�GG`V�g'7Y�Z
��@����C] �ψ�"\{��a����{zB�]�B}$�[��INq���`Nyc�C�ʧ9��� E���P��*���]-���N����9��Ʀ%�O�>%KA�K�a��J��O����w6.��ٙ(7�x�g����<a X��+Q�8�=�d�*�}�f$��^8Ie���~7��4ђ��0<�=��]����W��q���Ѱ{�<����23A�YW��zsl�j�!�d�w�$~F�^����VQ7�*�%p�{>f�s�	��;@�n�kْ�>���0�M1UWdj|���ˎ�V�g|�-P�p�+{"g��2+��r:g�Aw�Z.�o�+� 1/�xw��ȁs	�3�L��ڜ�#D�S�&�-0*Ag�il�eG��TJ���4)R������*!&s�,�[8ʧ@џ֖�Z�rMy��~6�����2�$im��)�݈�G�v���^�7z�P��:�U��b_2W�!��p�Q[�g\gC�?iA���:��	[�u�R]	��%ʔ0��wl���QJZ�Tޯ3vSLa�"�q_j�)�8��H��Q��7��jw�7#^������|ݩ=+}��@��+h��[��\�k��7�x=q���� P�c����uta�_�B�%����,<`�>5�Nl�����}��\�{4�T��_~����R\������_�����X5�<�1(���~,q8���rF)�E�C�+ �s=-��Ӈkׯzʢ�K��r���m��xr�����=T������)4\Ul/��{BȻ���t�8��Bi<�_)0+z�V��3���B`[?_��7��Q246��[��@H������（=HU�`r�Cw��ԣ�Y}�����7CѾ5Q�/���MMd}#���1�j��c6^X�T\��7+�u�ۏ��B�,�$���"�n{p��7��2� �aA��`�cg�)�L�T_����>~��Qe�Շ�qZ���#.�zEb��c#!�8jf�hȰ�`+�b3S�f]?�r�m�
٢�1d�{#�8��ʜ�	O��RP�� ,n��+���u`�J���r�U���9'�+0���H=F������^�~E���%A(�`1ª�'��g�H�2�#vɿ����LvO%m_��������(׍]�����#�i��Ϝ`
���"����q�C����%�{�&��	���]<������!k�A>Cy���b��A?+�L��_9ܿF��H=�kǣ�u���C�nN��ۺ^���	�;��i�P���9tɗ����L�0�L^��꫃,W?|{S�s6�s�f����Jۭ��Xqk�(�x7�g ��)�]�⏒���T{�������:G.�aF�F���{G-,Y�
�wĈI�b��lDi��\)w�����qs�W,�^�����%q�(�A�قE\LI�sF>�� �I5U� �NI?�h�� �V`FAF���_\��#�Tߛ�nOeg��dU�Bq�.#d,r��0���Ҷ�ysb��V`�kg�yHD8���l��"��cJ��p��ʕ��a\����:2C>�Bl1�ㅞH�4�q\�C��3��~�*��ހȶ���,�������i�1mp��r��Y��`�=D��VD�s��Y ��@�B��e#6-�����Ţy���mW!D
�X��|�b����� K>�Uq'N�
v$2��&�Q3�Xڈ�ōm^� �T�9��3�!�dm���`���Mx2s������P�zn���������#$�L��)��0S��;璜��eUI�N=��i����lW��M��}O��v]� ���1R��5�U�u:���A!���F mͩ���D���Oȑ\yzV�>�L��[u��������j��N�/�b��
��+�$�_�>5U��)�h�U�zŊ-
�*�z�h���W�W� 6�@�i�IZ�v>��5��Ҕ����	���ر�i�0��cxz�x'��o�&�#7�)��e	%��hlv��[}�_�T��j��uT
Y<णWAlҚ'v/�+��@�t����*�Occt���!�҇�;$Efݛys�ۚ��A��j�-`�A�g����D�j�����z8;��"�÷���v\��z�Q2�������"�MX*9�:wע����aa�X7m��d&���?�`>d&ձ���8�^e1��Z��x
$N�3�}�Z�"����gV�����&��J���(%�6N��e���uc�3��S��@d�M�`=�|������/�Bۗh��߽P�a�Q��a]���s!"wO��� KK��ϣG^���DO�|��fc���Z��w&�Hu���q�bW�ĺ�����&��Dzi��$	VF6˿��Nw� �j�_R�|�#B�=��k\r�UA����=۹R�р!����J�c�N�.�e�B͝2",a���̙�)�x�P�+cZC��H��\<�;��U���{F-��֬:���u`�B��q��\5��70k+����3�}��%�����&m�?�ߞ�j��(���^�d�+(�vi��l�1H��M�?\�Յ��E�t����#�F
���(��M�؀n�.T$�I���z��^��p\ �IE�4�;δ+o��ʲ��xW��y�Zi��Xk��e�"�i��߫:�2l<������I���3�W�kOZ�R�#�0U��M�[a?͵�N��~�b(?&�%�� �Y�������\��&�Ӳ�N���~o�	�u)ϋY`�-T��Fox$*[���R��&���3
g�*�����q�X�~~��ĂCe��?��J}G��E_}��F��1/)���9�O��g���H����Je4�ה��a�C��DM�EO�,h����2S�5��p�i��CXC�7; bg��(^|�.�~'G�)]�OrJw��Q�X9�����iq�������[<1[�*�����XG��G���ש��?m^9Y\�KYH�H/e"(� 8����P����oC���y�ę�e����Yo��b=�؁<�C<i7���f���JTrakʳO;=ynڈ�@~9	[!?���Z/�1K�k(5f�C��k[xƜ�s�nK�w�ߚwDoK��o<��z��RZ��y;���2?c�\�:!�0h}�iF�������a�L\R� @�P��W8����Q�/L�a�_E�o�p{��`|C0��hn�x�^�K�H�q_��Po�\з�֌��(��B#{��� 7��q<�|��w�tT��J��G��Y%OW��

G�05�U�ώ���O����ZM�q�K*v��%l)��f��*h�ϝ��;b	q*�IƆUD���>bɎol��{J�5`�Ű�Cz@V �u#��Q��פ��I�G�{�H&' ����L�����"�k�%w.M`o�b�}���!D@ioIv.(dJE�z����N|
㜊3�
��~/��UB�ڰ��v�)���9�"�E��.[ۓ���E'un�~Od��5���!d�������u`�jU ��U5� d��}�M��h�V:j��}��0R�m���x�c���ɨ��ЃQn��Hw�ގ3��Q̈́\�XzpV� ث<Q��~�0� (�Cn�xՁ��U�����V�E��Ss�=G;�����읷�&$��)�M��ş�(^/���g��.�����d�>W��A��z]�߲���N %�;��K��PcT	�(��,
7"��~�
�K�tj?~S����Q�p�顺���Ef��9V^�:�Vl5��0I�i���a�I�Kt�:U��ޞ�&����)%P��9���( �O��
�v��<�悇��MR���ɶ�-��-�����.o?��!he�
�()�+�ۊz69��N{A�6761�A����P����u��xNP���NU�1�괈w�����3*5��dɥ<~�EDC�vJ]���.`��ۤC*t��<�\x粦�o��6���p��J"L�F�,����je\>�g�s񦘆��U�>Kj(��{o�����-9U���!"�B��	U�4Ik"A�L� A(�}l�r�4Mf\�L�~��ⶕ�^B�������޾}'�Ԏ�}�ÿڶX�[�C�\��V���+��N��x �.�**��r!��&P�'�Kb�,��*%3>I������(Epp�������Iܮ���]�y9��]�C�R��qY2���y�}M>v�'��D��<��)�y�f��r��5�	�=���BG]��J�ߣ�� Rn���%xCaTs�ւ�<ǰ"��>P��"��9$�!̭@V其0k1�[^��±�d��B�ǚ9�qN��w��x_Z�`N]��`�zZ��4��D�����_��1u�
5o9&�'F��ӠG#�����Σ�����ED�j!ZLh��d;�ݕ٠�k^w'�^��8�Q�p��Za�T���x�44�yfjm�/�b�I����ł5��!�!cjjW*�~���7�Z� ��ܲ,qYdu��a8����В������=&�N&ˊx���^3�k��)�{���2)	)���U�y���+��:a��HP���Ov2��fW�� �x@ :�sީp�ǝ��A�hKi
v�v����������-A������	���Cf�%��'���s���A��t����H��g�]y���?"	�E��ŧ^���
z2���k{�>&������4���K ���*Cm�x�P#�c?�l�q�@��Jy���������'!�&�"S�z�g�y��Mf��ͪ�z��(t�ʝ@�$�,��X�O�Nc���N�ƠB�F%X�����SNW:�x���u8�IB�m˾�O��;s�H����V��u�|��Fr��#ߤqw�<̤���tº.�֛7���PC�o��	�\K$~烹0��J0q��~��� ��>J�ء(Ia���t�:4JJ�[|ҟ�Y�����Ks��[E�.x#� J�~���U])��`ҍ`����Ug�P��HL~�L��H�Lr\����9>8��5[p�p�)�РT?��к ���=���X��TH�$���!JV"Z��T ��]�H��"�� ���	ձ"yo,U�������Y�����3�(b��h�-��'w9��+)�6�)�KN��1%��t���^�i�����(F�����4DxCDT>�01qZ���hlP�;Ed]��~� ��+��ݭ����O�B����sb|������t����b0���3[�t�pL֨ŅT���wS����,�lǰ��ݏ��4����*9�V�}�F�IW�6�,�p�P��6�/C�Q��ekɈB�*�$����؞Au���F���Mk�B����\k���-K�Q�R)�諾ͯMu��LG:�2g��q[l~�Y`%v\v�
槆�H�t�\�)�$2�I���j�cA�R���x�����w��E�-��y2jm����:�Uu.�~Kc��F��b�BǐVg�)>QU�u��M�s�z�͋���4�Y���>%�}�$�T��Qlb��� E�7��?x:���X�i}C��Ō�C�$��@�xϤß�u�)��<D�=��� ��fs���,}(�f�&1��o�:a�R�8���Bu��c�~js�(s+���U�"�_�3d`��"�O�������|~*�x�E��t�[sZ�\,H�6�Ob<0���ob��\t�t�����j1;��*#��N�}��D����ϰ}�α�d��_����y�H���녞���:ǐk�Wj���M���T-���KH�I��8k�֑��P'���A����!^��:aǔoʄ����̗dX�P�;񩾵��,��Gہx"V��ή�u�`���`�Z����ޒ�ZY���HhT]�u �����c�B���5a%N5����5o(t?�y��H���.F�O(�H���17�A��6�~�&�Io�("�l�Q���$ﲅІ��1���Т���TyL��B��PC�;%Hۈ(p��r��	PP��I�h�}�ݭ6�a��1+�E�7{�Oi�D�;��x��8�{ �E$��\5͍��`�^�bn$���իI��fF���n��}��|hnz2�;x�/���f����}49io����X|�׳��D�R�p8�����)r{z�f:Z]���B�\ښ�F>��L~~ �Z4ލI+:���l� �f�6��I��c��*��tϠ���x�K�@6rS#Tճ�WF�����um�p�|��s![��L�T�^*�Qc>��lҪ�Uˁ��"h�;�<������s���U�u�yC�9 5�E1� 9\y�Ā ������܆,9">��<Z�����I��Z�~�GA�9�ĭ��~����g�Põ�2{z�X|��������{~��d���T<:�9#M��4m�Q�׳L������R�� �f��OuF�7�D�袖`�L��TJ���ZV{n`v���P�����]�+k�\�~;�MYqJ���(T~��D�(��O��&˨�_���sfHyT!�V!C�v�r��T���#���4(�l�$do�嫽k�;�#��̶���E]g��IO!��s@u��h?��Z�PSn�Riy�^pu?�~�a��/"9UZ)�����Ԃ����߳^6P���J���(v.��i���̫19Rin\��miV�q0��W8G<sr���� ���Q9NHa�fE���d�h��o����ϭ�E�ye�6��Q�r0V�{������G�S�� �c9�@�:��`C���G��b؞	|xq�O�[���|����,�m_�_-�)g���}���[����������iy�]�g(<dS�_��Uk8�R�Z7���$D�v���Bg���SΗ��sTy�<��$�/�a�����,�g(閲�w���t�}�����n5`;�r9���7HN�]�r�LYU�����9+(��!����ij^�'�e��{�.cZ�P�4�����\W��_Wg���C(�e�j���+�k����$��QN��Qд���_(Y,�t¨�O.�!���^Q��m�B5�Y-�������胤Õ����eV�'F�PFOm������}|�עs)W��H���	n��id�W��]b��!ڑ��/��J��	��ku�2j�b��z?��z��J1*��̢��/I����>��=��K�0�s\�T��v�h��u�N�}Y��M�������Z}#�����H�46Sk5Z���w�D��[^wX�t�J�},�G�Xiӓg:�<H$m�]���b��Wr��X�-�*o��+8�����w3+È4�]+�ک���v�����2��C��1���r��/%���'ع2�!�Vn��mj����<B�����U�w�~쥵q����Y��H�KC��YYq�(����Q�V�鲭Ɂ{���b{-?�� q���Ɔ a���h�t3�G��#U�qh��Ա�5�������>q��\�����,���ՆXG(�\�]*���P��І㟕�P|/A�jX}���<��k�+��߂��p6�@i9!���gZ�t5]CN:t���! ��&Ɣ�K7��li�Uf��at�G����W��9���@i��%��4ͽ-C<Y�P(��pL�=uq����C�=j;���)P�S	2�6N>���j�{�(�=ݥƫ���;�[�~E��V4s8�,�ڠyK=�٦�I`޾ۺ�M��m~=��q�Wڠ �3@� d�/h��%�$ phYZ�[hzgܜ�G�����-D�" 