��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ�������nu�-&(��v��.���j����fl
�Z�i��a�7�����}D��4�!3�51��la�%���0x�SzE�ڙ�Ngh����f�~)Ρ%^�R}�L+���y�%�8sf�� ���b/�R�@1�@5�ω#+��3��Ӯ;�6ȃ�`Xa����$�/�+{�$V=<m� �Y������DJ�(�Y�_�Ѱ��|��e��閯�ksY^�'�w��~�Q��۵��&�B�
��v���3�q�@�"��zK�z�l.8V"��E��\��I�]*W.	��G�E�2WIH�-9U��vb��ՠ��kG7��S�ђ�Sv��y���a�ո�����KW�DEU.u~�6Gwh'�\�nL.��;���Fϰ�ca��SF��3��0�yG􆅉HqR�=w�X�%���j9�r�����HC|���#OŤ�T@g��⡌f�Xդ��׋��c|H�����+��R*�L_����r�����1A��L��Q�%���@�$6!�e�\� �PQ�\��Z�H\�8�^y[��H��4|g�57xy�v�a�L@���>�l��pŨM���Iݲ�r���^\�RM&C� �����>ٵ�p�ZL����)L!�H�K�[�m>9�̓�g	K!�+a�F�m4���R"O^�>���eG���jR���V���z	硞Ih��l���͘�0 «n�u��ʇ�p�%�_1?5臟�*�H\�h�j\�]�'�A|P���$�#�hAȂ]��:�:�� O���ݾ�`��;�n6�|�T����fi%\�G�3��QsX%8�2��J�?\�'�w���MU)b?<�Q�E{��7�:�Q���a�U�~�d�Jd�2�рn���M����J��������B�d�w~��|"����9�I�Q��<�a�pa:q�O�û��7������j�Y��|���q��H�����fiÞ��M�7�G�w����SH��9`2I�Pٚ/��čr��c���~�I[:���Nk	�W�`��ާ����Oi''���3�Ճ�=�t��\��t��}���d��$d 3�_����X�E�Ǚ�(�H�j2����\_��lz�y��`ut�@-7��VTu}�����Ї�����F�yR�t%�e*q���6��L�������AJ!�}���
�I�c�|ϣ��1�ȸ�i������E߁x�:�#�Y��uv��U��f��"�%��^L�y��0lj�y��������K|�^|7\�	g�k��Xu0�o����#����ʭ��$�ʏ��yU)/�,xݡ��K�Yf-��CHP�ɦ�RU�(l��{m:����ِ�Z��a%�9�L�߬2*�(�l���x�Ļ7��*�;�w���6��cp�Q�:��ο���}�h�-�  ��0P��#:��9������3W�׭M�[��s����G���n��.Ֆ�����p����V>뷜Ek�٠OV�$3Q�\ʋ���ڰ.�����lhs��+xaj��L~VjZ�:��A��U�_3�T�u)��g�$Y��܍p2��,m�A#����h۱���D�/�ِރA�/�V:�x�A ��y�-�-`�fZ�$i�}��t=[ə !��Ջ]��J��o��|n�*Q|��z��#'��8��H}e��C8+]kZEuສ*^@8�*��CW�/� W���MM�6^۪��pOe+��Y7k�x�G�3$�W|��k|	/� ���^1�����]Џ+��ݹ�$���"�U[�S�U���&2�r�!M#g��Pf�T�V���x1?�G_�^Q/M���4ƾd�4�"FL�k��/��n[L�ɔ5�[/�0��ۮ�;Ӏ�7-�Y��<:���)���)v%�gE��1QmP�����禆�`"W��"��s���ꀢ���"Tz�7�ζ1�zi2x5�TQ��+�X�# hw٤Do�`o��I���w-U$a��������V�����X�,�ݼ!�	�cQ��:���|�Zxf��w�n*C�>���7�N���X�_�Q�ڱ��O�j�`�v!?�� ��Z	�*V���	Z��~¬l�Ǣ�y��{R������〣��EǊu"�bH�����D�` �׳�$��UDh���ĸ���|Z�]҅�$KV�@����#V8�U������	�%1�y�k�u؋��:Wϵf��m��x�KB�&��3�/p�x����Z5
$؍�����WM�*��*����y�ؿ���?4��� %��j��M���?����
(p3���{M wt��mM�tv6��؍ם��1_mS�b��/D�����]�H�;�����\z�	�z�W�,!J/�wr%L�wF��O�s�j1ҥ �0��$�-��+2�s�� ?��iy�ʮAb��(R�bT6``�s��U�-zA��=ǉ{��_���������浪K09Ť����B��Q�bF�
�U�-��"�e,�p\Tܓ�w��d	V# x� �J�N�@_��Պ^�}
��(�%}�o�|�Pg
L���6�6��hc#�~�����,���E��7�s��]z�[Mv���Ŵ�J�7�|u#�F�,�����?%W.smn�E��X��A!�V�P�CfʃlR��<}Cx�׋@�av��bvmt_���4z���Jү�{�W��[�l��5�]8b��
L���n���{,�vBNҍ����k�\1q�jD�n)QVYia����F���r��q��/�|d�*U�xͱ*9do�f�o�{���[�vxM���Q!
uWhC�4�0����u�w	��L��Zs�@W��7{Y�V}\+��ȯ*Z���hb]��;�v����aﰮ�Ed�M$��h������&������kā�����I{�b�hS2�H�3]ݮZmɈB�������*�n���:��E���x$�Af߲�Ğ��|F%dn~>櫕�S�|*����V����������t��q�"6%UFGd��f�T�w�,\V��dMxYJ�ع��4��֝�:�ҩu�l�ݠv�Q&�0"�����C`'��s\�zЀ��#n���=�h�tM���Kݫ*�$��CD�-o4�v 랫[�$@)u$�
�O�C��p��%��KnsaN�幮[zF,����)c�=f��<�GAsQK�1nR"{6��b{̙��Q��rP�	���F���X�Ƌ�ǅ�;e�a-�:y��)
��q��'����%�����ϖ��Yըf�g��/3�-�W��g#�|�дĄ�<�1V;9.D�m����
�<E��A�W��g�Y�ɯ���i��͆%�z�N�'�����p���Գ@&��ɕ�0q�~}:��,ڱA�4u��tĐ�������}8������O��� V�2� k�)s�,>�i'�T.r}�Amz2��y3�Y>������ׯt*���^`m�򴲩�y5�����l� ]ΔJ%QrB ��w����ay�d_ΰi���Q�R�����!�6�M�50�ls]��ش��og��y�j�w�e��|FW~�������6�!����/9A+�� �7����s�f�Q��?�y�ѱ}v@�N���s*�,|�U}P��:�T �94i�FhiO�a`�`H�t�BĽM�.�#�����0g�d����9�޳�ba�rUO��>��)g��C�?�	���JB@�e��;��J��v�PW���z\��AӪ�/*}��.5��qk*B`^��VO��L0���
��B��u$L@������{BЇ�W�U"�B��ʨ�;�r�tXtJ�6�O�ͤ�"4SKW�We����``�L�@Mi�f\�C�����v��;�C'NW3 ��K	GTi��uP�e���^ඖY�P_Zͥ��B��oy��YK������v�2x񤰥�M��?���5_c����:$��7�L���P�*Kʇy���`�x0q6��`ay/#14���,�6��`�����T�CH�V
��&�n�����P��<��B�Ɗ,���y[��EU��'>}Df,mV2+����M^����"�4xHar�[�y�)D����j6۽��s"����$���R�Q��L�D�0�k��������k8��X����`���(���	�`�ь���-{+,�;M��-�kV�m?�/���Ê^$<)I��i0��e��)V��49,�����n?}��tٵtg&I�����q�y0��ub#*OĊxw������92s]����.��)>�⚵��N�Uy����]�w�'P�aE�|G���!X�wg��BZ���GQ9��H8���R#��c��>�w`W�5�T������?N
ў9� 5z�0���߇&�i�*T���?ʪX�����!�oa�97��ܭ�aL�8�tɟLl�n�%i�L������Ұ��P�D�k�Tu�)H_a�΂��,���a��G�9���G�@z��Mڞ����%"����&`:��GŅo�r�M�����#k���w�n���.�m�������&+�̭�-w}t�\�D1k?c���-��"�H��x�5\A��m�5O��UY��̸�,�{v_�+jU�ܦ�|��dhI�x��K�x'��;����Vn�QR)=���;?��g���bd���~��OM���~_��u���	�|�q��}��
��B�^56��Nm�l��9ٚ1���֐5�7|G��\�5�)�N��ZXҳ7�n^z�d:�5�*�X��X�E�mŉ*
9N���=&|]�G��G������U-y��I��X��R��O�������BT�Ka�׋�(K�<��ꖴ�?
0J�?M;7���=�'��PG�3I�́2w�{��Ԅ��#yX�9w�L��l�m7���H��wN|^��A_��I���F��B��Zp9����E�T�U���!=o���n2���C�������O�D�{�f�]��|3��k��1��B�g-�ꄓ�Y:C�r�8G�-Q�L"M6�e�"�&wk92�H�g�p8�q�� XI;a���Y�ii������ ��T��|G>����|s��OG�O�3NN��
~vY�SZ%\�τ���|(�v~(1u�XO�[�K�k=��	��/���S'��C�v���F�j~ Q�v�	��\a ��ׂ��ҹp;_IԒ��(E����];�6������k����>n��M4��SL�� �F�Th��m|C��;�� ����vR(�ڜ�3��/+e�L@A'̒+��b`��J�{��?�9�7�P��M;����
��]�*'����7�Q�e�$�D�,�c�o����c�`o����*([�C����[@9�$��*fmf؈�f�5n��ai6��=?e�H�&��vl�z�w�xv��G�I�>��#]N��Gў�9���vv��d#|��ie��.D�
L"KZ=�G�NFCR@H�m�Sr˙�#X��G���f�R/�����An?�F��#��u��iY�s�o��UJc/Z����Hs�.n�e��6*��5����e(�Na��T�
#lOa�V{����t�d4p/�:He|O��~�mV3��5��9%q,cU�晇�vGmpG��9ȥ���є;�ձe��SUZ�^�s� �ٝ��`�y*�)��ۼ&� �h�2�U}�3��ʊ���sK)�V���Π�I
�D�G0���Ӆ�2u1�TYI�!��0Q�_� 16�)^����6�,�v;ME$P# �}���ɛ}�L[��T+����
Ͷ�����!#5��e+���OhJZBZ�;_n�B�4y��ƙ]B-̡��i�aF<���cyذؕ? ��"�Fq��t�/Cu��cE�v`��рb{�h.�F�8o|�P�$_����Fa�hˬ�.��G钰n,!���|'i��1����r�N/q5�����\+\#|0v�6�hn 4�~����Mn��_��A��t��r6�d��C�ȏ�~�2�L�,��������~��c��]�i���!#46��J��Wխ�V=]˰Q��N޽S0uv�Q
��ۖ��8� M{Yؘ�x�e����s�uov���Bד-�����={3#��{�V�9�I��ۋۮ���#�Dfo�o��i�Y�;y
,��jj�8]**�\�_��M���Hp�4�S�p� ��ie%)�`�=܏lV(��K)d�!�����b�]�N�ȇ�2���9��kBcZI�G�a>']���6'���&���0E��p/~G��6+>v�s�4-�x�A�12ޮw���C��[<�3�ֿEx:��ۂ��<47ÊCi'�ia60����}�R+^��F����B5�þ��{-��/��D��c�4hw��E�^�@괺��q���dz�_fƁ�3�KRX@���?�}��7�~g?u�x,@�2�D�AɺwX�E�C!m��k65�p(z�����l4�r0��}T��n�<�A�i�WK�s�V�hA�vt�AՏM��ͽ�G�J,qYS+�뫫ݮ<T�%V�W�2��B���vh	��>�f�K����* v�O����� ut,^8��[ �C怦(-:���}䛌gg6pY�p&����C��f2
({����<y�	��Ȑ�@aO��V՟8ޗ���˛�ިQ_��(���"���������Q�>�|Qr�Ф�R�b|O�"���y�"��PF�(P��YP�W�d<u.j�d��J N��tn[������
L��u���$�r���Y����Ψ������:�}����S����p�UhR�k9�����.�r�:CW:�\Z}}���}G��2_[n�k�!i����tV�I�O�xS�U��vJpu ��c7)sfg;�b�>ۍX-�^���{��>�0����!]H��!M��Q�iC;-���\Q�~s�S�	M΄@4��"�YS�	�
�ĸ��E`m����S��57e{��	��H;"���m�\!E�$s�(6�*A���ix���u��E{�fu\�f�;I��":��X�6_�U�:�BYƐ���$���,\*�cр_���'"iJ����U����ѮЂX��.����kr��
����8!�İ3��^}P�	`�[Y2��NI�{�Nk��J?��*(B�X��e�$(A�0�#����Z�κ�{PR�,�q�6#����d(�#�}�ÂВ����@���nt%�����`��/w�J17�2F���y�:7ge>8���皿���Ѷ"��-�^X�o�j�"Ȝ�SG{S���h��V�pT���u��ю*�.'�r?&ڷoŎk��;^�D�Bh|P�!�eeT%-%���R!���~L.7ܻ�\��8�"�U��;�%�6S'p-{ʿi,�M�S2eLA?� ofp����i�k&�?��,��� �Kڙ��5\$���[A�0 <�a\��&��hs�k�m��z����[�ګ'������e�%���-�|�:�ZrE��)�0d��D��w�}5e�o�¼<������_0�l�K�յ��C�dǮ} �夸��)��m��OqG�Ӂ+	w�p?�5*�����fm�pL�N6�!�w����0���B_LX��]�w��T2,gH?%x԰�[�Q��.�_{w	Bt��չ�HZ�0��vzy����5"fAG=�>X�����N�K�g��䫹I���Y?��Z<�}� 226�(ݻܙ�k��/�Z�-�TEl�s4=��lE�M�[whb/����ќ
+�D4�r��z~�s>�׮.]��:7� ��3���ӡ����g��]QЬ���F�
�`���7�?�{�&#���Ji�R$bF���8Mp��P�������LpF��y��h��̝��v��e�[����5 c>YY�D�c����;��v�:~���^����V���D���`��U��n�i'8�(Pϝ��J+e,�]���]gM��ii��y7nmf���A��j(���"�_^:�=o���O�Wa�87���J迼gW�j���B`E�&����M�[����A�J9ki�	c{{ %x�hk_��V����ݎo��>����8��.CE[�t?
�ǀ�ܾhʠa�l�B`�`I�d2�k9U5g��X�G��l��/��Y\�k�y�Y&."-��X��sTJ��Ŕ��]�q�Z|���������u�o�Wn�oJ�t�
%k�p}v��<�r#��o�ey'oq�gj�Bj�3�f�-=|�������YX���$�B��zB���=;�ف6=syD�I^�$'_w/����r�Oy�p��c��|�l�r����*�+���{־�>�)�����q�1_fG`'Uߘ��m�\I-"�"��l��\7�u dEF�!V~��� �gh�j���Wц���f�z�7ٱt�|����=,��<�L�U<h�_�e[	F�(�v�zGu_dSX��=ib�e`��=�w��=P!�N�oWѭm��9����B�Ǆ�`|�\��2Gb囹t����`ח��:��B�/��m�q?��s0N��K���Y��Qy�W �Z"��Q�ϩ���K��Qau>��C`�e����w��W�RB,�U�ե��
�<�����r�L!��GF��d�v<�H��(gN���L��O���e��C�y�Mw�'��k��p�O�SdT�G�T��}8\Fӻz�j�Й�4&ܩ�!A���.ݖnm����9�p�&a���o���'�%D,�:���l�j��"Y2\o{7��Q`̈́�F�-�
<�A���-$�<��������L���[�6W�O:�;���`�@]�4�X�}��I}����8�jr	y<���X��
�X�>�Ҳ��/��`����_�=���
�����MT��6"�n��R���lFy_�;�y���{��M�L܎�ϟ��Ԧ~$�0�zTa,�N-���+.�i�k���d�Tj2����=X���ra���v\��e�2�T��ٟ+���(���� X������ǻ�����J���u�>+�_
c3ϋ���{ým���f�����m��Y�z*�ެ��x�y�V>��U^�����\��D-�JY<�����t��%�?���ͪlcR�����쮷�d$�7t��%�O�4�C�~�xd����̤(
��"��F��=?eդܺ��d"�4N����;��Փ �ϡK�j����~�63C��S	�qk� ��G����+�;��k�.n���O|���c���M]���2Y��Ŭ�����{����*^TvC�q��C�<ĥ�s�w�����=���=88�v�ed����%틟H2Ϟ���7��2�iSG�cc���ߠ�_9#�g���ǜ�L���c:iɺϩ�r�v�8��]�������3m�EoY&,�����Z� 3�|m�Z��Uǯ_�z�ؙ"IlR��$h"`B��� ���Z;�*�(u�7�k��P2�����A?'ui�ר�M�㢐,k{̇�ow�T~+@cm�V]��p�dUJ�u�*�f	N�1 ��n9�0�o�������p�V:U�����&'j4�'�Sn3Oz��]��ߵel�G��MY6:�6�K%H���oH���=sv*XE�c��[����oz�i��r q�g07
r�w(D���~��G��M���i��ًx������|�|!�#�sw�����t�Ͷ��ps?��iX>��7j3dv@��8t7��j7��I�5K�����4Is�s� "�iR엕P����IH�
Q(Ҩ��2��;���G�E9��L�2Vk�V�^��6㧕�¨˽Z���v��̮��/S����1�~Ӄ���r�w�HT��^�슻K�x%�+�%�A�;�*����,Ԃ�� &;98=��h��'&n��C�;j=F(�7���� ��|�d�����&�����,������T�+?�H�ؔݟ��S�䧅��#�Fi�Dަ�%���#4��"&�O*���`Y�j�k ��4��g7s�Ț��3;N,�8pl5Zy�V��ȄY�#{��Ǉ���hiخѾ
���#j�>4�J�2��@'��0	�S���%O-�v�O#�_��������(�K={wC%�@�poK:��I`SXb��e=��{�e��P���kE �-1��J��f��w���!2�Y�OlJg�;�D^\ˢ��-�����v䄉�y�B�r�9�_��O�'p
c�u�ɍo`+_h�V�]c��u�B-x��cc���H�!����x ͜��@�v
w�B��qu��2��q��<�M.ٶ�R/�TAi��:9�O���蟧m�Gh=b��K�U�8~0�5,Q�9Zi��;�w�G�d�zs	�k6�R���o�oA��߯F��%�&-6�������3�&��Z��-�T�nA�' �(�@׶m@��0����$�� 8��HՋCpa ,���6=tL����f����a�P pq�}���joY~�kg���jw`�Fk�`�3�"�ӝ���K�
�G|�-t6n���׭��]�޼��c�6Ў��XfHϝ�si�4��ڟ�d�JYGbT�������I���~D,�e@��=�"�I:���~�q�3�N��~+;�maB�z��nS���<;I���y%R�	�l�n8�
����՝B��뫴��x�@ �3$t{x5ﷳj��[o��@,5�l �#FUm�ӚOo��.��6����x�bbצ=��A,t��D��� ���=D6�t�|�v�[hYz�F�x���5,{�@ޝ�q�-�գ�^U�)�fGp�+�̺ƶ�ʮ��,����[�<�,�O�I4.I���U�~lh�3-&�+����tE��u�sm�4�� ��[_��y�1�Ch>������q�f����O򪋴�|�7��UƺO��緤��J.��U�k yg7:b�ThX