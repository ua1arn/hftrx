��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�Ck%���-Yڙ}VmCt�"=��Kv����7T'���b�ұ��mڧ��ދmϩ%��=��R��}���\����N{��]�+,����a��@*x��ƅ���"�f�{<��g��F�cpE�)sX�m�k6���P���vW���Ͳ��&�].��x�	�+�bMM4 =P���ΜO�x��?�̍���`'~8��N姃���?�qt�`�5�;>�(k����p&���Cݪ�Z�<}x��	��aC��TG��¤�j�FxH^2B:ڙ��渉N2������r�&�K?������ܺ�Н�]�7�7�j�F
Q,È���+%�`��ةQ�:��b�����$���!�h�Y!���B.s6.R�J|`j�<9h���-Q�{�U4���t�:=�(3�m���3�X�R���{����2�t�7��e�ۗ�����f�c��Ӭ�K}�ｔ�MV���@>ihM�0�I�3�{OUj��
����@�{v�����Z��H��%?X�~!��؎u+02-C\#�c�5���@�s7�^��I�_q���=���U��Jw��
�	���'tVp�-�)G��$LƶhnH�Ra��[��%'�Okˤ�&�U�]T ��@?O���Hyͅ �$���b��Ca�vo��Y4���\��	\ TS����+	�6�b+���]H����0����>��'d�����<��BU�ģl�L<������񟲥o�n�l����l9�����vQܐy(3΅�4�|�w����S�B'�����By�&
���QCD���j񒢥~4&�o�����a��:��ܤA�#U���D�h�_8��P����� ���ѿf�V�UN$��KJ��sCZw�2�s����N~X }���T�9qb���¨�}��γ�I���d��;.PY��y#"��n�  BEaf��瞧U�o<�h�GU�}X��R�ֈ� ��T������٥�z���< A7�1���Av�rkZl����Y�C=>�ݮ�s�w0������V�O�ؤءْ�ulT`Q|�T�ȃ!i^����2LI:��B`�F�o{s�g�:�hf���
]W�8f�)��<����>��l�U:�uIK2�@�t���V1+�C<�0�>"V{"s��Ј��OBsD���F�����j���H9��a�.E��=�n�q�f^b.-�V�#yJ74������tX`N�쬸M��se��Y�?�;'��,���E#4e�⭎�T���u��0s�d$~܇�D8�D ��X�_X�)M�4T����B�������+�w�]s��{��S��m8������ +d@- 7���}.�.aX��k;�m��M�fa��Þ��2�E*�����=��4���B㟸SXg'Vh���`YLύ�z�;�ۯy�	0��hT����-4�w�'+#�S??�g�J���.�T ��Q���s3��E�Z��vW+X�ɥT�h�+��&<r�������a�a��棈~_�'YN�a��d���թ��6Y�4i0�EV�H��n.��)�K�p'a3 :��B��<N��*&������Hڵ|��I�8!�V���!����,�\���q�E��C�]��ު��Ņiò���7�-�"N�3�a��?�=��4 �`i�i�C��υ 7,�9;$r�4��`�<���&�v����Uw-�Y�i��`x��Q ���E��ΝWЄ���x{\�D��?��P���K/_�5U�7����gq�m<+�} g������<f$�cl4U��D��h7���m�H��T@�����n��WD���"r�������M�%��b�ԋˤ[E�0&1оA/�/7�mҮ	F����"��c����庂`_��DT.��?3�~���L����S��<E�WRUlCq�\ü��J�f	�G_*�a6���q�k�ϟ}�D����T��^���a38�ujEQ�C����^����ū�.`�+��ؾg83R۽c����~=1qq9*���+��O����l�lz-�!�3�~�9��2����}�ɂop`�U�z��S?����U���h#�M��L-�1���U|�~�^UE�աk�󐭭�k����������5[�_S��L�\��Ũ�V����Z��h�}���TmH4�J7삞�Ou߉�}@�S/0Q0�7�u�����(�H*q��W
P���+�sk|m��Rg38�4��s{T-ku�~R<��������H.<�]�0���k�D0�Ilܾ�(��{E���t�U�F�ը"{~�*�6B���:�8�/��q�����f�+�wV��)7;��L#���u����<������^�=-Z�T"e��f,�E���Ȼ�dWq�46 � X)e ��Q������@!�fK�����~q��7rG����н�y*�����ḃkԭ ����{��u�% K�8KP�,MjB8�:N����.���wbl����2�^轅����])0��iWhg�����޷�\2xX'��G-�V�Q�sgѵlXQ#�b��0Y�nր��#@��]c��z�Ұ�fQY m�����P�j�8p���RE�*��}�sZ�RJ��i]1x��N�������܍t�˘(�8Fʦ�^��m������Y�ɺ|�#=ӱA�����V��v�4i���/��%p�;��-�A�Ӌ�5�$`Ȇ>���\bQgr}P^8-�.X�a��t ��/��q9�ּ�G��nt��%��:�#V�<Un\%W�)AN��&��	�]#?+�ʹU�T��u��t���_(��<��]3)�sp��U:�Q�	Q� 0@[!G�ZQ��gM׈$kA�c|60U�v�D����Gq�:�a��H|���='#�SX=L�/7u�ȌC8Wi�T�ȭCk� �H�����λ�Q�i�r�GڛU#闣�}&��B~US|�R��d���G�)�u�T&q��13~ǭ_��)���9;i�z���9��ؖ1 F����eLs���p#�����2�#T��r�9|�0�D
� ���s��U�C��,��9�C��5Z8}��[%2���)�?����*��F�w�i�r�h�[��!bp���,���-�������������������霩`�+���������|�Cb�\,a�?����~�{;�ؕ����/��ƕ�Q���^!�o������Dv���-a���L�.�麬���P���j�)%�z��ӡ#6���s<C�tM.�,�VkH6���Gc�����ץn݋0sj�k���!�'�:����wg���tq���WF�ix��ɞ�fJ�����7Z�n�3'[���
q'Ī䍫2�&3�Jmkm��g�V��@��҄�����I�Ͳ�)Q�౯�(��MEv���n����5�΢�i�,��1�\��ŐJk(�c}���w�w�?{)���?�f4`�KR���َ�L^	���C��ŷ�\�'�@��-�c�k�Wĳ�ro��,'�w��"�]|Y�?���G�rFg�P%Ǉ���S^ϣ��5/����>U)T'��)O����#K��B�;�f}�^�K�$2�	�S3���Þ� ����Ä��;U' ���BPCpJÁ����e��pEe�����(�����q��8���Tu@q��@���q�[IG� ��E�@���`=�;lB��L��|�-m>��ح��TҌ�Rw��"bG���˗o�/Hk 0��6$�:��S�ͥ|a����<x��nU�t*�.+�3���#T,�T�bZ6 ��U�D�[d�_��:�C����LV��Ix7r��`��ҝӛm�h��*�e� PK�Т��xH�a����9T�?�53��A8J�}ȷ�ÈP�����A��PL���2.< &
�p��3��Ek���fSR���������8�$�*���Mk�j ~Y-P:\�>���$��K�P�f�5ȓ%|��-�P��Ft������M����L�j\3�.̮�a��^�A���K�䫈�V�n�]:�MfX9]��A�(�S���+����'�c��_e%R�<��A�F�W{Wa&�6�$�{D��� *�}�R����,Mgx$��X����qI�.���ž���e�M8�ﾮwѼp�
)����&�M�nP��:�~�T7c���F��J22�l�����](�v��O�6�)I-^#�	Զ?�f��+.��
�����'D���W�L�̗4e��-	g�� `�a*ʶ� ��a~����t���&^���j�`�#8�ӟ�nLt�w���u��23Z�� [�BV��L��|�h��N��Z�w\��.��cZ�1@���=�����9�+:�*��	�#��O�����EP��H�),�PӖ�.�<�j*��^��8D�=�8&�2���1k�}�Æ;^ܩ�-��dV�*����5\�%�>��g{I�#o��ˣ s�ɫ��#�t��,i�Fؔ���:=�?(�=��'k��6�Yi
+�W.W�/L�ɸ�BoxS`<ڙ�������GvL@ےXG-��kIǱ����5r+_�K�.��Z�y_���M�p��df�>S�2�%���RDD����]C^�Ʊ�3��B�T0�q��
��b�a��K���J8<�����+��3n_��Q�nqD��_��2!�����V-PB��F�3Bx\�쉸��A��+�
���k�,ܵ3��`�P���~~$t	we����>��r�ˀIm} �ݖ��Dmj\1݃�p�(���}���P���Z�ԙ�Pv"���mg�j����A�T���X��l�Rf�w����R�`�b!��N:��ŭW�Zޘ0���3��ɏ
��'�,ğ���}�0<C����x%���8�fw������F��\���4FJ�B�[��j)S���L(T�c,�D��0�f�{�zp1�I7(K%�Q��}:�����q��<���_�������UX�����q��a:|}���-zӧ�o�ͱ�zH��å��=�%���Y�	D4Ά�c�n�����Qs\M�+�x�,;��ֺS|B��>D�[+��"g;#?�D�=S��ȾR�|c�H�Y~�΂�=��.B���f�:���-�W?�=O���,�ď֑��~��w#�T$�/��x1��iP�l��oe�X㟏�i�^'h;@@�$x��d҂g�5w�	g-�!��JP�����. ��������Y��!�ߵ>��:bcz�b��'�͏Xl��@}��y�1, �8�GrԤ�����+�$�T��?�:1T	��f��f4&�����Vn?�:�)�o(N[�|%�R�W��O/(=�`s<�]�D�e��5)�?�e��Qx�m�D���N
J�_և�Ʋ���
�l佌����܍"�C:KvӼ���E\�1a�%��dc�l��N���O&r5z��HñR�3����^��Q�2���|�V�ù���=�7bL.�H¼~�������g��[��	��������-�k�셭�h,;b\PGB׍�R�R�kJ��a������ �%��,J��ߩ��j$�=ԋb2��j�z睛
������L�X~<d�WH�Mu�s&�%�{T����%��ǉ>��@���V:W)���d%�H�&us�)JS�q���O	�'�1��`��k���n��:���zV��	��u�z���cG��C�����c�*	G�w�>|���HS��]A��#s%��d�p��iC�T٢��{3�E	}��+�G?��u�#�U�n8]B�i�i^)p
��G�E%��>=D��m�O��!�VG�7q	�*��b22/�|����h��J�� ���K@��/�k4u�,vJ	!���}.��	� �������3H�&���G�".��ks�rf��/�H��������������^neE�?����)${�������7�D׮j�f���[����Ae�n���21,�~�i]v��/��ˮ⥗9�c�ˤq������.bL��7u�+W��/�w��S,�ϯ�"x�Y�cw�9M�|3}b��Ҏ��	�v2� V��؉��o)th��^�6�)��lƙ�p���`<K���j��_�/O+�M��n��^W�i>�Dp@]\���
[b�m�J���.��3���l3����C�v!��B��l�a0����S�:P����`�OQU��q��ʒ�����ɼm�3�_��� r5O^�����u&�1����|���R-���F���aȸGu�³9���;������%�����?v��9��E�$��}����������B���W��,���
������S�1k��EEK�*�O�%T]g~��|ż]5����u����H�>�*�X>f�VU�&��&bE���H�꩗�W�~k�z��+e��`*��m�,��Fx���U�
->]ߘ[>�x���Թ߁����I�\��pl��~7�5�uSgP��\.>��G�4͢�tc���s�y�+��AC�o(t��K�U&�����+�9�_b�~P�>�noW`�Ƒ.�[US�\��g���6͢y�Y�CV�t�<�1p{�t��_���n���n�z�,!G'ہ���F��l9�����ؚ8�*�e� ��<��_p�e$���o���{��rr��}(�p�q���D+�}Tk���^eG��RK&�~��)e�5����&�/��z��@R�.�~��\���_db��.�RGx#T9� ���Q���D�܆��ょ�t]Z��j��"@O�cdÄ5��ҙ��L��	T���3���o�k�q�7��%��͵��%K˿�8�6/��5j������}N.c�����s#�:�Ji��/s�ɇҨ���h�# 	9%Zy�	S������ybR޾�1t�H��j���t��rF���MC4�9�C~����s�!�E��B2@�[��F:n?Ψ��<�\<6��a2ʪ��\~ξ�,�p9&�����B˽�4r��T���{r<�LCԯ�U���������?$F�Jc�`yǙa�j�w�O����A����[��:T0�,��8W
��t����V T�<t����n��e�ü���G�Oځ�Ӟ���X����:NN�c2vK %r����DD��U�R�(Ҕ�7�&�85y��^�����Q�R��/=z�)�d����W��n���8��|��_n/7M��Ӓ!���0?�r��x�J_PL71�c��Nz����-���&!�9:�b�vI���=��%L�f\��b�M�ð�V��X�{�\/�IhX�5tW����O���iR���t�'�9=��a^��s�)}�ږPژ�,��L���k:�:烖���?�i�4]��=]�|bm�����X����j��Y�0���w�09�W�7�J��݀��}�˩K`�:ӁD�k��<��c< )���j�Wң��{�S��[!��l�H �l�4}���i;�d.؊����.,���/p8,:���H�<��R�>�.��atF��W��,�M�.[���t�A�W?O�C������</�$z���[(�>�b�Y���Q}^� �^��Wq%32f> �{�kbw��k��T4���.�f6�8H6��Uf���#�X�@<M�q���c����2���`�a�9��*jE�X�A���]�'Q���q�Y1�e{0I�mŔQ�7��o3Rmz���OA}�9�h��.U����M@�^í��j��G�"@�BcQā� ��;?�}b&�v3���:�B��b��+���zr�ӷ�cI��yۜʒ��h�Ԋ���4�єX�^w[Z`na��f�b� cB�M_ܑ%;�\֗A��TFڡ�����p�~�X=��taʫ��]�_�������9I�������v��!Ų(8����#��(5��b�����-_��׏i�x�;s���c����<��ȴ�;_�]�$OQ��{�Ȝ���4RJ��<�`�5���S��������3Z�*������MD�S}�v�T	��jJlG��S�Jb��Cr��>�6�'��GQ�l5�"�Tb��<f�c����յ���k�}u�+d�F2����z������8wCF#i�\�7Vg0@XN�2��Gm��^`�����V�?�_��&�,B��m!��δT�d�ɸm�R��L��:���W�f���:��'<�ւ]l:��������܄ Ǿ�0�˝ҍ z�K�_xp:�Q��{��T��J�@��ϲ'��NjT�`�ը!uY�/N�j5A6د7o�4A�d��Lҡ�Z�;�9~yF#��G�n�"�lj�$���RV� l�|>�Ko�e��
���,,����{�(�'d�c:�?۸e�I��	7���@B�tm��ڃJƐ���"X�>Y(6�ஔ�C�.~E'�qe)�oܢ�g;�������Au��ͺ�n��N�l[\	���n<���Q���Kg�X�3xh���hk�djM�y����G ���D{̝����Sǧ�K��3��{$DN�����@��'h �U��<���L���6��S4O�q�ze��XzH����V�_O�t���fk�^��.��5_�ver��/�-���oo���8Zڏ���wg�9�����<K_����]�����w_ �"w�K9k�� ����$.Iq�}";�m.]
o�ʺ1RfO0I�Y����� ^�[��-X�KG��x��X�?D;�&�e�7@��Oaw�ʼ��	���a~av=%W4H��f�'��(צO��X�r8.���Nb[H��!�� M�Y'!:7~~��!��(�	*4D\M�1�6}x����a�rߓ�n ��3���b���Ϯ�κ�o ��R�.��֝�J+��D�-�vV���w��䄫N{�UI�\���;Q���K	n-WX�4oQx����=|�P�|�	�p�X�]����B_�ܰ�Y��@���H��qV5*�?���t�Q�Ё�X��x�~?�b�[X�"��V���Q�Rar��X 5�m"4�Q���ʆb���A&3C,�;M��C�Z^̞PaZ<zţ���m�جH5�#�z���z �C_9������_�(J�s=62̚��7:H'*�PL��u�t�AG�r�X���� ,��r���i�XWP�Ng�
��� ��Ag ��l!�M}A+��ӎ�E=�I"?���O��7OH�k��:E\�d�t�L�f5pw���5��0�{��-���Y��	-ߘb	R�V��uo���"ҬD�c���w/}.�en����Y'�v5
��~J�$�Q�Ϣwdߑ=_�}�0�4p�u��u����2���>k�b+�����t �V�9rq<�Z;�<Ϭ�����¥�i���h��A��c[������7�>Q�g|���<�t4=�J���gvv]�$�-k[Ԓ�OJ箂<>�(�dcJ�o�FN���w�C���G�!R�$m�dZc�t�����UN��3,�T* �9�0�J=�k��I���7<{aG�ͭ���F_A� ���{K��[Bi�ʶ�M4�ވMqm�D��!j�,OQGn׳��B�{��8�y�0����Ҹ^�0�z1�	�>�e�ڇQx��ג���SeѦP�~�8�m�j���AK�����T(�	Ųʙ�����@ґH������� �RT�K��ԍ�3��?�@�����֖��,i�Q�X76�`|j��"���H�3� v��3(z�q��Ս�x����+e�Y��
�`l,U]*�2�4��zq$��j������jơ^Tk,^�pޘ��%jv"K�ň�_$|��-j<ċ�~LM)�y�ak&>��^Ş��T���kȗ|�\�>-��*y_�T҂��RC��.�%����8)�DTǥw��&rw��r,�A�m	�uQ��m�6�)IF�+�f]M���)O�f�OE�� P�^�{���b=�k��r�:�U�5_xE���D߲�a�*��
P�V4s>�Y����@T-yd`����m�?z�T��J���xhP�RŠM�3�~�(�!P�Y@�~5�)J�Vd�w§���$�oJzW4OldN� ���D��+:�`��;��G�H��B�ʙ�C=*�$��@͘�����X~�7ܧ�����nY��x�X	�($
�[q�ǭ�xA�H������Ls�cӊ�_�f*����S�"@�lҏ\J�������������$��2c�n������Lh`Z	Y)
U[��7D��u�7�\4`��Q�6�IC]u����f����6�
%�T�x��ɩ�=�����P���d���	9�u�.��%�s0#�d�_����F.9�|�۽Mz{�ƸC��lz�7꽦�����T�Tk>�r>�#�w�)Gs���J��B7��"�Լ�q��dx�
o/b�]+T$��Ki��l�g�H��0hJ�+���k� ����1�>o���ٍ�e�H�j��j���'Mp�XBc�������8VEJ���p��m#.��[0<�6���+'�Ȃ���{��_z}�9�?�/v�-�m�rފa4�[-��2����]�z��0��{���{���c7��Zo�+��o��!}ǝ>-B��0�H���å�#�C�ʱi!�������tG��᝖.���EFiW��ut��g�h[�v.p��5&j	�A�C��Y������h����Ms:�M �Ʊ���k�
G�L���`	�����m��u�	���!�):e6���<�N�:�̨M
)��]�]D^�O�L����
���e���f�ԂR���4i�=��O-K~�f�!nHW�����A�� m����# ����ℒǱ�Dr�hx�x-X�U#��/"9=��f&�9���:y$�J� ��-,+m��y��o�&�$ �< XµPN&?t��C���6�s��q���Ҽ�1� �F\��(�7��(LA�ʈqG�J8u�T�}���x�?��~��RD�U���� ��rv��s/�څ�eJU�̍��h�㙯[i-d��G��u��G)NC���5����*h����z������a�{�Yx����ȨP���9�����9�)H�ɕh�~z�")$�E;=�"��B�Q�R�ʣ!��|�d��ug[艟^+!�Ӯ���w��|���oN���8G���R�탘�¡�^�IM�q�2�.� �N�G5��ן@,w���+����K(�{[�A�2~��{�I��d�C��"��?�ڦz�%��5#��g��v<�"g֣�vfq=��]�	]��.�vd��B�����M�_�8�P�jV"��b���W���-rqU�Ne�Z%�2��!	��x�Hc�)�������vI�h%D%0�m�GڀG�6r�-�?C�T���pb�Ğ��GV�1o�&<o8��e4���q��,J{�@���m+��2���\\FWp,�oy������5__�-�de°��/�Q��6����4��d�c�0��*�v]���]��`�U�Y��0�c^����5T
;MƬ����3VH-?Ap�:.�L;���r����3�H�7�?���������}3o���;��n�#����$�ʸQt�p�Z��"�3e��e���
G��L#�o9��F;l����OȨ=d����e�&V_I�j�/"Ѐ
�Ixh��K�X�p\�<�.�xY��a�G�wK�J�E�s��ui�Ԁؚ�7J��#�
�߬Ĵ���$Z�U�X��<�x� lq�n.K�N�d�y��� 0���&��[6�8����' �H�����##��c)b��GB���_5�H�5�������e��c�&.�'1�v�2z�4�O��U-,�W :�b�S���K��`��>��o���|������2p��:�BVb�N��b����p��b����;�}J5L*����_��I��R%�C�j���5醎t�0?j��j"�숮MQm���������;�`�_������G��\�W��Q�:ɽFq��V)h�:��o���e'tA�@��"��xn��b?�E�**��Y���;ڳ�{��:d&'�%�Zkw�*�Cg�Vq����5Xg�'<����#D��'3�oh�o�i�*
�h�L�~p���[�w�6����W�wJ�{�Y�����Ҡ
��V+����x=��t�.M?��6���Nޱ1D���O5�݆�c��y�v����y�uE��{���}��M+p��܀��g5���C����S���D�#g/�ӓ�?Ǎ�)	{G�`�d8�����sE N�e� �x>ɿ�NX�~��A�����	w�o�{���B�`�Q��Rr��?,����n���z��kvm_őR��9�K$�"Z0���n�����v�+�g�H_�Ɓ�i���*���K�(��RJ��f�pZa�W�L��Am�w  �>EB4���_�9����D5���0��=�:�zj��;3�e���J��"'���ぬg���/6��1��7�p+ͦ��w�OR�ֶ����1`_5s�!\��
��S����?p��&5O�ٻ�{Y,(l*;���҆�Kp<a�m�;c�Z5!����N�u�{� �<�<˳�
K�G�Yc:�%�eb�HՆ�1&�i��ue�W��F��qq�s��;�Һ��6i����r~l��)w@U���d�g���̐���j�}��nP�Ze*�x�X���F|����~��ǌ�w�a�L����A��/�@{_ AV�N�����FN���f�4S�j`!���<��\��0���]���/�z��)�M��~��f�v8��!4��
Ĕ6_z���ǰ��$3v��_��~,/�|��ɒ�F�W���i��v��+י���xQU��|�w�c)�yZ�$vK�kN�=�Oc��n��+��xO)����d�����spm� ώ�K���]Ĝ΄K	�=�Hi�"����������x���
� �#�1&�,�6�b#�V�B����Y�����9K��[��*!~\;�o������#%�vU�ȧ��v��x~��2��ġ�c	e�\ZQ��H`贴�e`��|��P̈́E���W΅vLF�Q����[SQ,B�$��u����, �t��D��{/��}3+P�q�	��kHn:�C��R�b�@G�����,���;
<�`�<�k1���s	�4R,Dvx�AEб�Ȉ� .�ø5v�H��I�9:�E�E"�-����j�z<"�����%,���K�3Wʵ��D^B����$;U0P�ó�;�q���e��Ɲ��Fv!���(6_�Ċԯ�7�s�̫h�m�sȚ���C v�`Y~#ܯ�0X�a���_s	(�����Y�(��k�(5�Aph��*��>)��W���>���$+Ԙ_���S���颂���W�8��{�	�5{�t�.�h�q�PkH1�#�	0	#��|q����A�`�K��8>�I4j'bk4����w�w�w1���'�k7�Pr�n���ɪ�j1�m-z��A���Ǳ*Ć>�#d��¢ɭw�h���!�F"��YDuZ�~!�!�RK�RS%�>�V��?��4�au�Ç�L��HO�9h6���m���>7h>��Xu�	��y�Р2Yҏ��q�85�,8���2?}�_��g��Y58y�3H~��-��thiHc�g��v	п�7J�g�m��Oq&D����S� �{(i���2M!��X��v��L�t�����َq��`!<��~˅�O$�'z�CC�bF�R�}���=�� �7�R�*"�`��TDD��hR�(x�\���	��F:ٟA�����,����������ʠW���	P0"�D�Ҡ��\Uk��J� �FS/]M�m�|�U�6��0�"�U��5��corD'�oӑ�|���_m���ʹ�֘�>�;Uy;ӯǚ	ϖ�ܣӊ�j?l;��� �4�~kB#��3��vpG#wE���Q���l���Q�Y\�Li����)rx�/2I��4p�T���葡j�_1��zi�����S��_?�	�|�"A��@�ɫ��+c/@��s�i=8Ά7�OZi����@�h2|Y1��׽��r<���8�IQ���,�s
�s�4l/�I�j�yX�1;����; �(��KD��UsEsO!$�#⨓�];��g���"�Z"f�P��bU"����?�h@7��0�2�M��E6E��O �:���k�?:A�1�Z?�(�x�u�B9�^�\�]~f1�c>lԫ���Z3A��)ê��c�E��_jO�%{ ��R7��l���4K����x$���ň��ĝr�U��]�b�ښ6��u]mPL~+���P8DA��q��U���co�����:t[Lr�>)9\�J�x(x�J��jɪ�p����b.p���#��2�I�U/	����7]��,\�߼���R��ytt�;���[�7s��PϠ�$7����H\�ab��x���gV�W|����X)Lv.B��I��p=���.;; �!A�x`����	�#�I���'�!C¦��K!܁�c�o.%,�^�d��J~��w\��Dm@� ,�ɤ����`���8����r0��m 8��hp="����q�Y0��Kf4P���a�[CV��l�1��fn��t�I��t�՝��1�6�/Ⱦ����S58,;�hex�Qܐ��(�0�g�l�i>�H�iefV��M������P٧X�,�Wg�~`{#�7��|�*��L,�['��-w������y�@�xa�^���v9�-C�Қ����W׈t����9��4�sFc��W���K����9��8d 9��m���'T[U�e2�I_(�ֳ��@iw�C�u���0�D��̈a�ˈ�V�^2�ݮ���3�I�.�
~01|�W`�F�Ǩ}���K�Ww�(Dg6O�h��4	��=�&�ZS�m&�[�:ziJ��1u�ET�Gv:i�x�W�rc��(��P��su;x���D����tH�e����`t��}��L�m5B�%�{���/�u���f�Ut�Kiʘ����L��Dڐ$��?�c�Lg"��+�΅�8V��}~s�l�#���U}�^�˱^�+��)1��~>1n�bo:b�Ԝv��C��K��څB�:�Y��~}�rW���A<u�)aط7SM8��3K������$���4��sM��(1֍]y�j �x�^��T:.�`�$쪛\i�~rt	d�W}	��z�@^\��G(�^���B�'����4��Dy��:�#{���������I�(̅�3y�@נ7���.��\4Z9�^e��,F��O.��6yP�5N/)͑.�Щd�@_ӓ=:ʬ�bo�ݘFj�⸥i)���=l�vÃ7�?��;��ۀ?)-��ѿ`5�mX���5���e��wc9�"%�E5�F�Gg�a	@�Tw�V�"E�-_R
ӟu"o	.�i)o���6��y�b�����#I�F�FDʕƥ�˛Yۨ:l	
���0{aJ��e�C؀MS~*�-�0����ہ߯�\�Z,��w/L�i��İ\1�Ù~><�]�0�(ɞ�d�J
�;�������ޮ�3��dҘiZԘ%�SS�khi,��q�\`E��LXwb`4-1pl����&�Ti���|'=DG��;ÏNi�Ss�/�QP�S��J����%��N�k>�_#4"4�ɨ��`[���d��ljӚ�j���m��ZJ>7iۍ���TU>Zͺ�0�eX=h�HqLFIg5��2\5[�o2���Msl�E�Α]�PTbK�,Ox�|��m :3@�+v�z�°dT<�_��^�zT�s#_U kQ�e �'=2V)���j�ޖ�I��xl��!sD�	�f��Ad��.�`�V�Ip�I]�bA��K������-i�}P��}��	��GSJ����iK���E;�����l=�g�dbL� ;f��{��(Nl�V�"7Ғ�̡�����q6�Y�硱I�Fy����I����:��PPf#�G%x���ީ�:�D�R)i����&�k�-��R�H5N|����+�́�Ć�u���WA�t+�=�����Z� 0S@'�B�{���aY��]�D&�����"D�{�{�nA1��L �i%.��M����8�)1V�Q�fJ�ٙ'�1*!�&�՜ W���;~u�j��Z�Y�ə��qjR�m�������goK�A�f�+��F�!h�f��د+�|���ㅬPeF����+��VӨqf�}�s;�E\�Ա�1Zu�DM�����$�gI����D(n����6�hc
�U�h>���(I٣��έ1�e>�?��)>М��K6:$�:S�h���gQ8`�����e�T*]9�������e�6�O������C��+C-�cn�wN�����=�3ʝ�yA�VO���Z����Y������ ��U�'�
��4�f���E�<����]��������H�����B��j_j�ǔ�QR�t|=�aI�r�^~���al�0��om�	C:9i�v�h�\Z�tz�"����Įʇ�Z���З�)o_ᣄP��,H23O�>��g����2޳n�R���l��*����D��D���3[�~�4�eh몱O\��RU
�"����EZ��g��F�-�/ݺ��x^�����w�xk��������C���;���JC��%��B��KLBc,�$��-���<X�9��#b�����а߽!$�o;6!W|GΥ2궅�2P�+��@1ܕF�n �ӝ���*�79w��RDB����1��3_lCD��KχA_-Y>L�wU0�J|XS��4�?���������o]���J�¯x'�� U�"{�r��/��N,MD���b��'Y�T�kh�zʰ��\ύAum���n�x̻g��B�0�0����Hl}�0}̙��w�o5Yz�3���Ԅ��Ų�A��~���8AY<�r�+�w�����i�F�߻�3G��h�S�=�gp���k[�����:S����������,�,#���񵘀�a./k���E�܌��8���N���kL쓀s��"4�9�y��[�zҐ�FS3%����p���ő�d�}���s���W0A�<���>ſɠT���*��� �2[f>D����Ƃ�$x9�y���E�Y�f�1"DV��Oq���`�x���=��Rb�;o5	�b��J�jdG�,�FJI�i�Ի.;�P�7��Q�h��kSE��
*���F���|B������=�7x��3"�����u��4�������_��%�O	螨46	-��S~�$�=(p ��T쎳i�������Ҳ��Ǭ9��L;���Y��I���"2|e�9�����%��AJOI6��h]�?��P}t:���!>�EfU=�@�|��kho��L��Kz��Q;��-���1��\v��咽Z�	�&h�~��׭��K�*L�2���I	�j��r�������D:�k֣���٩��%���1�������|#ԃ�.UF����c֜����\��C�foʀ[ΔG�d�'VA$l�h4�׋����Q�τ3���ľ�Ϲ)��Z�2!��=>.Q�A�:\�����hy%xI�*=�F!�����w�K8 ��[4���$p~fD���i��(�ݒp�]��38MվL^�����w��M0E�6�.?�*��NÒj�݉Z�g�hn%��/t-�Q�K�B�G��"�`��enJ�]�w�]�\�-���ٻ�'�;�?c�ҝc��6��tk�{D��|��"�u@�~�D����I	�$��G�e�"V�X�ӧ4�?,˔�T~��D5=�f�"G1.|A�0m@����w��������s�S��H!�#YvVl9���%��g"��bj-ۆD5���*8�)��1U��v����h�޻U�W!,����q8�I
�����G3G�4�G���c<ݝ�����b�+|LM�'�"c=L_@�'N�Ք�� ��̥B*3��w�)�71����E�H����+ �|ec�f����\ñ�U`��5<[�W>��|���N9y�����`�!s��� �|�5p\#61$1�M0�	��D�%o�F��.�M;|<b�n�#o�h��;~n�n�zj>����hN_��N6��ȄPn�g����A8���<��6�<xtd��!d��Nn�  �0s��!�c�|;�D�r�� '����Hh�6����B�h��f�<����O���Ω��!Ek�o���i۲�W)]���TUoj��ߒ����H�YjX;ʃ�G�^|�%�ͣ�rE�����|�ۨ�U�|�T״��v�{���ި�x2w�#6���#��V����h���g>�oW3��٥#]����ÞaES��P2�������T%�ʼ��߻��[m'(�	��s�/�E��S5��W�0rD
�3�����x�mz���
,M�s��@n0�=/�K������b�]�G��ɣ{�B��q<����e$\A��y�%��>ق@�[[��#���f`��cȬ�w��LY��MVI�ȥ��;��1cOG�*���,��i'C��}�?��O1Զ&���=��mi!"O���dŦ��g��d�Z2��W��%�I۝����
n��5�p�O��-�l���d,́�b #9���z��
_G����� ��|�)8���
��mWM�=��Y�b@&�c�fW<(I}��S��O]�kO�{���|�K1� ���w�t�Jn�ʂb�Bz�~ I����;N�s��������B���+�����a�a�ޓ���>i��+pE�#���Ԝߙ|Ĥ*\<���L��d%��]&V*9\�)�-V���	��\H7n�7�	�HFZsH����q�w�&�7�khAtn�XC �b��("�����"6��q��U�����wp�#p�
2>;�׋jW5�=ǹ|���_)�⹋W]3�:�S�}ɫ\t��4�����x�-D��9-����~��_s�D`�B	��KS��ȮF��A N�B)�yӰ�Өٰ�<��T1��v�JAJ�i�L�7���i����/e�+�	�op"��}K@.-3m���'��3cd��ƥOn�V5�7��f�X7.�~*lՃG�p{K�#�r���BW��th��=R1 �ACpk|�;�hݥ��\���փ��<��_׽gZj��������X6�/ѧ�-�!'���38L�`��ʜ�v+ш� L[�C7�@8��w�i:i����a���j��:xb|�Zn�#���w��%�iZ�E�B�_�XF���D̖�֕�?��������8S ��x�{[<�<�]�!)K'�%�,*�d�`���J2�G� '
����׍J�5j(;���}�����<|zF&�v�+����uO·�~�6/a
X!]V�sm�=��0�}H�W�zUPR��<	5�>�ǖg�0,���s�������y�-�p�M
d��!��F!gq�a���֯���>ʧo�u�=���!Z��L�� ��,�/�N��)5�j��	4pC:�r�d��Cѣ4|��P?PIj���+e���k�*A��x��A�QV����;���	�j������`� ���9`�c�RLrY�A���]���w��\�t�]i
��T�'�2֕`?��另����OX5\�z��Z&����j��;��^b�h
?M`���-�o��)���X�Bq�����⬣n��#;`Q�Y�R�FY�)��2�f�t,*�4�Y�B����0����H�45�)�1��+ğXQ��B��F�j���]%WT� "溼��wd�5e_]!�y4;h�鈈�W��zs���9��S�����D������^7z���ۜ�O�@^�嵘w-����?
�Cl��v���{Z�`^�6��,�uGЁ��0�-ok�˄yA#~>oPCeO�#S���%Į�����r�"f��s���Lb��x���͘lD�
�bk�&�%؇� w����Q@�$V6(��5YeP�����i��$g���t���\+��β�ž0���z�g���alq4Y��[�[�s�ROV�,��E���1��!gkP8>��bE�T��4 /��j\��6�)�i�)Z�FUǰ����}����8��d	��χSIʙ�+��雲�}v�.`+����.)��|.rX����q��$�o=�|+�;I�DQ�T���$��.0�.9�S�C��,��̣�Ǉ�C1͂h�Q�nͩ�k�&��� :���A�A�lcn�-�=�-O#$�#�*=6�O���Ƚb6$sh�*i�ϗ����y�}����lg���_�PB��YO��ɬ�ۦ\]>+,}Ϡ~�R���nG�0�uW��ӆԩ�i{d�D6����WM¨��������̄�ɄfJK�A'�X&�I���B�}{
=G����ڢ����f��y�v���",3����"ӆ��p:m���O]3-F�C[UV��0���yx�m�J�����r�0BgM�1;��#c�(g��X����!�w8{)�&]��?�p�;�=�sr�C�����=�|Pi`�b,�qۄ��1|�;m�S!�� N��r�����@�J�ٝ~���u�������-����ՃDt\$Kf. ���:�iG�ڐ�^�j.�.�M�q �������Z�\+Q�0�qo�K�#
Y��ҽ���=��D��w�j��]����G@$T���,0Tv��ω)���B��z�mX=՞d�y���Q�#�Z�]�Ӣ�<
�y��8,M�Z,KcǊ�����+wvq�=���B�?
'��H�;�⒞ueN�|~��f9�*3�8O}����Z�n��VU֠�~�8�M<ݱO~׸���f�?7Q��x�+g��&F�6ށw��}Vq���)�=�<n�..�Qs�QN!7ٗ�uIM��>�j�\��ʼg���`Y��~�����	o3��o.GO��]��n4ҟ�˓�	ߝ����'����n5��! {��T�B�D�Ijo�)�C��~�і9��ft�g��U��9���M��b��o�<��𙩿�q߿rɰ`n�����)���;�9X��f�̑��~���%� �O��g����\+��S���6��$IȪ��n�>^w��`�hFv��]��ݺ*���AS�໠W��&/ϛ�X�Tf5B�5�14�t�ƕ ��- 	���5P<��@p��`L_|5h�*Z�){����z��]5概���7�b��ьL�`�r����A k,	_=AF�=6�S���i!� !�"|��~��
��m������|��s��E�C�� ���O�<Ұz4S�PM�#���\o&��,�x�"[gv�"WFG�z�m���!�Q���x��R����p�'��mx�2_����<.<@bVz�:2��wʬ��y��Edݜ8�V&���#�[�!������GS�
�t9�GK�F#�p��=�QR�ǎe�)�h[���>�>R�������J��7MIpA����s�k���UJ���JŦ2����=+-��oi����XQ$��\��4UE�-U�)&�c���\F�D�1�˽��,�{�Б�D�xR�P�D�dĦ�?�%5�Ip*���_,����9��c{⫩�M�^�e��w��q���V*Z�q�qE�,�4Ne�q�������x�e�8�r#Ԇ9��:eXߠ�S�^M����2=Y�,wh��X���͐�KS��t��b�l�D%�r=���Sp�3�E�����V�<9��\^��;`t?��=��mT��	��,p�{v{� �߿~.T�Ф� 0}~�SY�bV�{ߍ
�V���Fw�op|�
�����ۛ��.�&��#۾�<��ȯb\ �sS<c,��%�<�o	�x��uF�L������b������H$N�4W[ȧ>��ݔ=�d�K7j>xn�Ï[�08ZK�w����j4;��B	�P_{fz�*�|}^*m4�E��7�"AA����
��l�9������i��#k�y7�-�:����q���;-�a[S{�u�����
��c�g��"��,kҷĴn���T������i?o�~�@���T��Y��'���b������^C�l}�6uƩ��EW=i���(�=wmƗ��wccb�q�p��ڽ��ſ7�5
��1�&������v[ȿH�+������4�<v:I@&Y4�^돇p���=HrD`��$��m��G�/�-�/��PY.�>&���Չq�q�W޾��1b����rV�j2�����`��j�"t��\�fxBlt�H���� �e�pe�T��ׯ�ѫ�f@&� ���t��am������+u4]��-]N�'�2b8�r��o��$�A}�����H��P"JQ~v��[w2`���p5�KR1��'�(�w��8��*J��mߨ}�;Pl���}N�u���d��Iϩ���o�����ayG�v�]�F��:���7�A�rv�D��;^�^h� �����|�q497肮�o@��%D��9�\	V�/��Λ�t{��Y�Jx���e�N�S���:'�_�vw����Ӌ�s�ף�5MX)�廈�ȿc�Z:9���_�-x�4ġQU1S���lR�4�ck�%��x��4P`�ռ���/)�5>N�(��5=����&	��_i�K8��4�߳sZ&��_�?��B� �/o]��YH<���;��J
�~T%��)�
�EΡX�ǰ#/��Ȑ/:>�'IΫ�q�h�,9�����$ �<���i�\��A+z�LUӲ�)?Ǟ�>"�*��O�)��#6!�l������Y3h���1pp^��n�  7��&���`Q \�DX�D.R��Ӣ��{8	��{9i�`_��-�R�t���t������դ,�P:�,NS���%"`���<�����ѳ�����S��N k�J��Ѹf��^;�~�M4���4�R���)C���L�k��9/R+�b�?5]��G15y�x�m6� .OA�KY5�c(�*�^]�4��>�H�f1߫o������f��������� �ڱ]�%��`�ss�rY���ܓ��,����l�ZP#�F��C��S3��=�|+���>� [�-,����*�Μ6�8�`tė1M���A���D����	��y�M�aJ�U��	�F��%c,��nNy	 �����9�M��x�~��T;���.4�<#zbj���͟�E83+`#b%�恧��J�&���mb*���{A�w��zw��������(g����v�(í�Χ��A�D�����^��]c:%oUJ�XH��$�!ä��p��I�}J� �	�u�:�f���a���TtT!��#����cr���Q��m�.q�h��݈�%+(SĐ�=� �i_��f�BnPhC�;����+��d5�y���{���.�Z�@:<B|i�Q��>+�R�������������rLp��\S��K�����q�ÿ@�_������- �
�Z�䪵��ݩ�6�B)�*q������Yt,m��:O�Q~\A�bF�0#��,H.xo�ӆ���NOK�}��Ȼ]��i�E]�����#���T9Ҽ�d���
���/�(�v�d���|�����l|h�G�����������"R�V�,�{"D,^fʰG:^Y�i��5�%�H� R�V%v�A�����I͍�ZO$�s�
U�����K� ԋe�ZS\ã���ӂN���1��B$}̿3o��x�2O��_S�1��يBXq�m�Ӝ62}t�R%��.�����D�kS\�n�}�Q(_x"0�n��K�'�镢��X����u��ݐ/Rq�%�tA��Y~��R��I$j3:Q�Ȭ=�5c�R�HE7�^wh���D ��)��y\��Y�6k�抹��9{���c�$����}s楴�%޺j���P�/*�]���~�E)��,�j$�E?n/�഍æ=��A*7�QC9���$�"�B@U�$y|�����C9uQ�����]L__�RF�m r�(�>���V)���.��4a����!�əM����?�@���ױ�	�?�S@�˙M�����W�l�1g�t��H620�}��щܚ�5�@�3�lԾ9\hާ5FNJ<����㟝S�\QB'����1��i�^�����|5����(@&L�P��p�RG���V��^
�-���I��Z�جxO���~]Z��>���Vhk4��Piu�"t�ry@����0�ɿ�Xt�Hor��ĻXFS��ݷ#��V��>����4�i,�X�1,��O�(3��@0��[�6=��+!|E��9t���i��b�xT� �zw©&�ѻ�Sx�"�'��dk`�o�^�@++�aF_�羅�Z�㫀F�"��F�gLARi_�i��#G!f��^g�-���~�G1Тd^�8��F����@`��P�4���S�{2��a�6'��58:]�L
��f %:�tU�{��9P2'8>$i�t(��#y���@���E�8C�`�L80�.���a"E,���P}��{+��C0�� ��@����22}�Q;��.�0=xU�MZ���)��C�5|x�v��:�8t>vU�LkտV�q(u/��|���1��L�:/��_D	Ј �W����x��T�h9����h�q�����`tqד�G��ϰ������=0j>T�A�� �jc�R4U =k�b5k��V��׫X��p�����Q�?��g�Ps�-���O�B�b⽼/���|��L$iq"���v�cT�*jr=>�B�r@�J�UysQ�c�T�c�!��!�Y��=Ѐ���[�6׳��%z�S%~�F���`�1W�:EC��
�B����]�(���E�d?P,�gɧB��ґ㮞~�w
��W�����Bʡ��^�[�ӂ]��7�}�x2�r��e辂�0�K����0��ʙS��KܯqW]�]��AƋ��9�\ۯIB~ˊߦ{r�
o�뽛�(�$`͜7�2�Y8�,�&�o@���s�b�G���Ɍڗ���3���Sq�ޑsl�`r�i�Sj ��׈�(v'��]�2tKW,\�M�3���C���}*l;�s���p���Yj^�:)&J�C�I9FQ��"�)�b�+y�v%k���WY	gXh�������,5O��6�/������^ds���z�Q#v+*�_No���H�y�#)
q���F��{�������_�����|0�2F(F�Q.����7!=<��� 01Ż.��Q�
5U�D`Jķ˫�G�0WJ]rS�W��4� L��PIbz�Rq��R��r"��RDn�h��l<F����^Sc����!�ȍO_��BB��>�%�R�~���C�/`�j��B��"m돸��f��;`��,�{����$���a?R���#������|8�]G������=�,�\e��U;�5�[��d9��/��_��V��'<���_ǢP��Q�C��q��A2p(�j���\a�9}�]T��?���?TK`����E�wЖ����4mW�_f�����\RP�je� S��a��L{�B�UF:����K�槮�7ع�&�>C;X�Ӆ�&R�Ax�s��[��B˄�Z����w���j9�K=��&��~
"\y)@s���_ �������ԗ[�a,L<6��䡌�^i�H]=��O�W��Q�SS-�����`�z"�΢@0������s���Im�-�ն)x7�7�UI2{IIB���Lmٙ��M��ϝ���3c��֗�U/b������]jAe�n,C՛�y)M�+{�)��;r�i]׆š_z����~?��
b�ֲ�i'/�rE�!nb"z�-}��I�N��H�Bm�
)������k���H:v��|�ݐ�1*.�W0��w� ��uy�Y;Ҡ�M��Ș��*�@c���ѻ��Y���	�|u?����ow�戫0���V�KE^�[��\)��EG�ݟ�
��),y7�<e8�J����	��C2�Md����"�i�@{d��.��Z�lY����������Z�ݕ�ʱ� ��{0�9�b:B_½�>P�[�c�r�2��=" j�G��6��p��u#��q��O��	)~k�a�q�=2�(�2>8w/�J��p��!�n9�E�1aD�>����-�-F�17΍1+v���saTj_i�����%s��yG��P�����U$�Or���,����A�#��
_��
�KR��;��A,�z�۱挃3f��b����`"���-�QiЇ���w��l���m�>�������m]���I�w�K�SK I� p�KzϨ���6�F[��Y��jIg���>
�J�^�QP-\���=,�L6�*]��tI�C�!B��DZ�u66h�d�`�X/��uJl6�-�ДПr<�<]�⣯~۴4Vj}z���M�b���XM�i�\�;�0Zf�g�Є�DPaz���a�m�.pN$<^I }�S���aYZY<z/ޘ�"B��z
�6�ͷ��Q�6�??ѯ��I��gU�H��.�ŝ�+�nm3@§Ϩk͒�q�M�i��ueK��c�C��dǈ�-J��j ��y~BAP�g�,0��o\���"ۘ�&���(���ۍ��x��pA�bx jے�e�L���06��U�1`�n�D�4D�� ��H}�8O}����ؠՔ�Zے�a!�T>Y�U��ܔq�>���� �gO� m�=oX��(z�k�C���&�J��7���2��^i�g��ڇ`���Weq�z��|W/�q�J�[�I,fc�ߠ�z`�bܦ����7�-���/y��-7+p]�oFԱ����d�e8���]}����G7��UABW� �~\KY2����`|�5²��f�&����Հ���ol���luW���5l��42<�֊L\9{"��_���_�x����������*�ӣҽ�G�y>�i�/��yIX�üVX�x�nds����!ZBE��e��t�qJ-�WW8����e�K�������A�Ez�&������ⷮ��'��ϴDUS`������M^��������^�l��&��o��N�=߉�k��;�3)>gG�zNX�2��)>l��H^��c=�C�Z<�A�Iˋ�c��+ҟ�������rji��SrB?�%�0�g�~��{�Ku���B����J�#"p�k?���Џ����m���O���7��.W���48`B��cR����v���'6�Q��oI*�(�}��d�<��ׅ�}�\���ρ����py'�� /�B[e��a,�Z�o|���|�hǓ��J6�,P�V�?�=����E�R�����fadrG-� �U�fN��S ��+R�7�+�/�7�1��q���]���sC�o��|��UD'�Ū�C��~g�T43욀v��5Y���غ��2����3C�d��	4��\�X�Ex��	d5'�s �����s)�G�����^��^��b�,�,'/�	�ct����}kk�Zu-��ES����6�&��U(fO����p�c���Wp������ˏ��k3���aE�	[B�{^�Dld34�[܀X�����BxI>�E��F����̈��������5Ad+f魫�ZQ��HZ��y��k��8�����|��L�1�
N���ӵ���!�H�Q�hT����%�a��4�B<��1y� �lD{�w0 �+��eAn�Q�d$�8v�A�|ǳ��Ώ9�Z\�똪�3X�Z;R�Mj��sg��j�259����t�o<%�y�:l�9َ�Ź)f�'7�D���!S�א���ƚ�<!b	<}�A����;�n�<�M�Qy��)��,ӱ�����-�Wx�V���5�����m$p�[~�'��9]þj�7�����'��l'�C/�J��L��.Ú6?�P�]������W�\��C��7��ƿO�Pq`�t���q'
�(�S�B�Ψ��b^	�	��QA�m�DuNʍ���&��:LXDZ �4��S� Ԯ-���}�kJ,\S� ,r��m?�5!1��Y��Y��fm���*�����iج��ب�]2-kd��K����p7[R�M��s��%eΘ�џړ�/>�Q#|>�.,]�ѓH��#�Fۥ�g���^P���C�w?�O����^�qUe6�5D���e�<|
?�`�&7X.��,��Sf'u�K�����$FQ��Bz�W��C'��_��G�Xn Q�<@�#����둕�x���W�L� {�5=�����=~��z�*A��!�~R����}}Ogtk�[�|�����J�<�3�EĦ
�V�F�:��D'�y�r�Ӿ�i�BU �o���cx���;OQ�i�x� �wC߹�T��-�3O��G6�o�}KC�5v�b�{�@I)`��1��8Ō��my�4�V���_7�ߠ�*��+��.뮃���Uw��=X�u�yU�D�Gz~RhA��w����BL��g�
c�{6��bp��]2�%U+���"���g��w���Y�~�{/�'w|) �L��_���c�qs�A�m�eۃKr�M_j���ă�4nl��uk"��ti)U�Y��ujcM�	��iU_��}�0�u.u恝� V�2�5�%�#��o�;Ԝ�+큍oז��|凌��j21�8.���@VerF^A�}�Z����٢+]M��-�u�r�>0bdbď~!44��1�N2��R���,�.����Z��̓[n�+�v�ğ����� ����k���7X��i��H����Ӥ ���l�
[�F5����i�\4�hN�h���������D,x�Z�"��ං����(-N+�����n�7���9����3	z���8h��~buCp
��-�֣J6���K��������
��"uN��>L�(�|Ԩ3�JRDLF/��~>�q��7�y�ʇ+-{���OS��/�1H9c�s��Z��k�%�N��(�&)7���G�p�Z�uE��3���/�xbb�K�1�rz�	@o1L���fT�'���ę�V�[If��M�X]pM��c�{�������*�d�y!"d.e��+�ۮ�]��d�z�<Xx�����Rc�S_��nF�ٍ��� �v�GeHZ����� �3�/�#���8���^g-���{za���{]��o>
�CH������_R�i_�$s�W�3��B��9�����nz�<Ҙf�����3��r7��i7����D[�d����&�`rx!=u���6��28���7Q-q��f��ھ��zr�ޭ����9�
-E�J>gUF)m@�=;�l��[�EiA� C�:U�$� Ό2Q �	<��N^����zSLC����K�-����Q-�пڟ�L�8�R�}Ў:���P;Z�h�BG;�a�N����\ya��v�T���
8Snb��R2&:���g:/v����&v��O�����N�U���@!yEjB���%���K<� 7����O�� n�T��iGF�F�H�- ��Bi�3g�A.~��-t+88h��e��*�V!����W����}�{P#�7-���\M���~h �����fD.�D�m�|f�6�A�M9�`oB80�<W��R���#����5�l[T�lfq����Fn�6���W�������Is��� �=�ވe)��(��t5$�+O���u`�[}<���ݹ�%*�U����䐹�r���5��Ƹ�F��&$����UG�(A��O5|(���.t��K�MXG�E@�Il&�dD=mk�î�Zhr7pb 8�Q�>�a����wQ���?��by#.J��j��8�#m����y{ D�Vf\~ ����.7H�o	j���T&�V�e`�m�>�|2�6�&<�|x�({���ͼ���U*pߖcj���vrD�c"k5?�B~�wBxi�$t��l��6&�CR���f��MP��+L���)R��0�.'}��w>����j��6닣�=|�JC�[B�Ms%~H��Y�DH�z�b$�M�\�Y���`�H3��G:��e8aU1��-�P�U�"��<����֛-l���xK����{���BRr6Nh�	�07.��H�M��(�02�ެS8cl�{Q���Ë�x���}��~���ԅ~���^�b8��l[f�eԔ�����$-q���*7�B+��@�B��ڮFP�wZl�e�*w�ػ$��8"E��
bV��+�=�ڵ;�8����f��k؈�����S�n@�%=�"rJ��_����{1?ЃӐ!<���7q��7I���`Jo.�1�����5*�V4�8S-.�q��Z����� � ��b�7�޼�c����tV��#��A-�Re�Dގ��4�����~�}i�e	H��!��`Fq��r|�}MJ�j3O�'�$V�xeL�.(T2]�V�B`H�h4���U��}��4�����."�AY�g�S�C����֔�m��Đ��#c�Xޒ��uN��$��=�)�HOn�[���˚�8�Ѫg(P'��)��z*N��Td~M�yL��4vR��D�(���| 4&��w�7	�|�{���wW��_�1��B���i���'�*�>\�7�ï̦%�0a�|�v�P���IJ	pTMr
Ny�;��Y8l�t}b/l��A/D���?((km���;��R¥�Yt�>��*�d��C��`�H_IO��(t���`�����!"����?�L�;_4�/��9�;}����R�A�h�U���i���1\����5G+lTP������h�
��Mh�.��V]n��M�p��l�?Ɨ�!��O�m�fc:ˣE��麘��s9���Ͽ�^�Y��b��0'��^о��kSi[�og�kf�T>�Bov�!�fdl�.�b�n�`��� �pD1X��lY�qk�E�!��:#��Jnh^��z�#v�b��P=_������;L3�ɏ�.7m�5:��xbMŠ}����pҹ�Y�F�����B%��m��}�	/��j��+a}3�ʍ�3{���r���+@Qq@�X~Iy�^y�@�K��������t!�%�L���o��������t��,
*���܀�=�Z6ǉ����7Ԅ�6���� a�hV�pQͩӢ^��e���E��O��i3�+� 7e�-�M���Di륄݀�xj��2_�����X��Z�����?���M��i������� F�M��|�S�H�WU�ʠH �忤o�W��G	U~�F0�d�jk�z��hp��c
�Ʋ��9��c��#��*�D��ҙV
�a72'<2ߜE9'�����ԌQ�Db L�j�6,]��ӨN^H����eqx����+9�ix'V8x���(IC�'MNW������B,=�+�&zò�w�2�R��]{F��q(�ά;��}� &iS���8��
��[	s�8�&	�;�D(fה�>1h�d����⳨�V�����Kct2��t5��x	��P��wt{�G=���"���|h������U==����y#����/HO��=#}?�(���v/���~�q�Z��!i� 8"�?n3���2Jd�U���Ɨ����=�t��k�P�n��T�����4�<�F�ND}/��3����S�����O����GP4�T+��l2���X��w	CFd\�)0��2��kn�,��r n��?��Z�GsoS7�N5O�(-U4uN��	��Vk���̝����g����Ci��B
x��9FĢ�XRu�W���m�r+#4���;I��B���ۺՇ�.�:��;�`\���d�y�H��*��P|:���]nLƬ��r *a�\݀n��*:NFV�hH���@��ԙ���K8��Ͼf��u/��W8�H'f�_�$;�n��!�Xͽ_Pe����͒s�C�Ќ`����q������N��)Qd�-���ض�;(��3;�"t�p�*�؁��L��TIS����?j��� U�y���a�[��ݖ�ԏ��-[���d��s\!>]�%���֧���ܹIN� ����ƨT�6���>*_m��G=�"&C- �3���G;/�S;T�N�d�3�7�"�0g�I%�M}�~��r����h�bF<��ʓ��C�ȴp��ޗ���ȭ[��Z/v�G۪�|�מxq�L�h�z�x~Lw�>7�%&v�v?h�\�+�������i�U�8����3����F�p�c��)����f�I�V�7�j:3w���h�M�D��nj���P��$��A���e�����T�_-˂_���:��m�Z��8$��\�.��?���>����z#�S�V	'x�7�ڭ�EԶ�l���$T��1bRS��`��=��㰗�'QX��$ :z�jh@�B�3;��FQ�)re�c��} ��Fؐ�hgs9$����D���j�B08�?�١�����*R:������}F;��>]W#�6�*#�¤{?�5�1�2M����; !\cyP0��;ǰ�>{�6q,r�6����[�=U6R@a�6&�Xk"�%��m�� �hZ	���o�s��l$;if���HJ΄��45��q��n���֘��B�g�Њz[ᵔ��<�t*��>��b���a��9�e`�#tG���5�
h��q��v�mZ�1���B���pǤ2���R�~e�I}8h2��8�b[��9n��`�nKy>%��@�.Q�e�'
	FD����R����ǸjKѶwN�pX�g���y8�"���^�^+�6c��Y��'�(xg�{E'{�0�"�dM�yB3�S�*oQ�t;
q�z�okw�!H?����ա�{GM��ؙ���A�X��O����LE��Xb�w3�~��v#"ӡ-kg3��胢ǼcQ��e���װ71�'z�0��C����#mWlw
ڛ���A��+ݛ(6K`d�h� m��(���J�lʬ;T�0*����#�Ky@�T�<��4��x��7p�9U��wU�E��2�����{!Sky
��w#���)�e 5�*	�J�:�[u����Z'Q�7���e(y�;�k��<Ki'��&�ԕߓ�5�,v.k��(��a��E2���nVԔ����3�8�T�>�u̜7N���L4�E0��svj��O���Uc��(�jxb��gQ@Ygа����E4��.�ʆ$��*�����=�8��o%�f�#�-��r�	!��uu�N66ޒ�{<o�i�� j��q�B؅�3z1��"�����%~�Z�*`g��0�i�:d�4ҙm��8jmq@��jS�8�L8],o:'b��9#&�p�՚\?�4��i��<�����"�k��hy�p���Y�h)�����ߎct�-{_h��dHPk:�`����~eF�@���4��hh�Q)�6��&��1�����n¢gtM��m%���[�Q�
�	�t�+MB;�~�R�|�*t�ՌU��벃P�\����!l�����i�=���!��@��BI'b�(XKl�4�h���%:䗊����,|j�OtxA	���WkQ�$05��C��,��N�:Q;��{�C�6�]M��gwo:�q��"Vx	ʽ,=!�����?ʄ�>[��H�C��Ԛ�G7F5N���)TE��Bs\l�o��h�ް-)p8�0�أ�/3�> ����Vҵo.��,߂� ��W�l�	Y����������cQ�4�X�{�/Z1(�w]�g����U�ݙ��v*�6�N�'EK澙T�z��@�<��'�:��zH�ͫDbz���W�t8�o%@q�d�Gb9k���u�F�k����x�=��Z�S=ɚ��6j��"��	�7��C����h��B����5��h��.낮E'�YL�2D��H��a���oK<�\��T04�?������0�%�Ri��8���m���}�H�~�4iF�s�^��es���z��[��Jq.����W�c�����
�����:�tWm��t[a�3�#���#�8��"�_�b��bQ�[:cӲQ���w�.9g��R�	J)���`xj�|��3lQϭH88�B��0�������	Z�X�1 g��Q���p�p�o�ӣ8����S��)��ݼ]aNU9t@1y;�ٙ���q�_�X�ۃ����W<�����l�r�6����`�=\L�w�U�1A��A�����H �D�s]u���n�� @p�5qX�X��A(X��8U�a�w���O�Xs� e�טI���B���cc�@�� &m��73�W@�|όk"/�b� ƥ�L��z=�܀q<�!�$	#�4� 2-`��-{�r?e��Kx��k�g�-�ߝ�㗤�|��)�>��{��c��yf�%W0GӲ�1M��z��W�y��d�'eZ���.�ܪ��4~�~�
��˳�@�`cT��/��A<��\r��wU�Ӡ�,a@�f�`�o�ŷܟ�ضFZ�a>h�4�[/��{d���'�s�X<g�{9�M �!ct8m��} �-�n0T5ؒp��D�TwI��σk�%6/��	婅.iH;�Oh�`�7���/G��F]р>?ک�h�墍5S^�1�����]ϷR��1n ��}�e�AH+)�xZFeC�//�=���`�Kנ�s�j����pf�yi�C�㔥�ħ�C�8�i��~����C���������B| & �C�'����\̸@R����&�6�A�~��j��M����o�m��8�[�+��{<s��]b
���K.K�B�3��ɞ�C+�O�t8��'=f�w���k�\����F����eX�P-diٙ_��|��<1Y�U��^�-�l�@S����45Sb?F�=�v �f��|�g8�udb�J��4���n�x�C����
JY���-�!��	��5$9DdnR���ޯ�>̷(A(^�����������;��b�a�f08�D]����}|�U+���?����֤�Rݳ�"��4w�w)�Ưo�.�?�!������ |x��Nf�%��������F�h^�~2k���ǖI!f�H�U�U����_�X`���1^G�fh
.V���@?��@��h5�^�:��r�~_6�5Khq8���ϓ��1�t&�eQ<yw���O{�IO�k��K��Q��`��rl(�t	�Z���>���P\qya	���joYP�jd� ������ݪ�a���姞���K%Kf���%��o�p�?M�v��2�2�p�SL%5�,�Fria�5�3i�@�d"N
����:�0��/��ĉ�en����a�[���a�\��.�a��[�j�t�w���J��U�a���7<{z�_)��/ň55w��s�E\��dg��K�W�h��F������3�\����3�@�N�{({�"��X�ٕ�@N�ň[���4�Nlz/T���z;m�>?/E�r^.�a*�5�X!�Z�Xe�,[U4�\�	L�M�8����T �j���[�4r%��CU�K��n�Uԑƹqd�o5�%	��k�c�&�7����$?%����QL0BLB��H HK��v���a�^�'���4���<�9U�T!�b�hw��[���bS2g2��6@t����z�&|�*O�	����H�'K��<�`_1*�6X�  ��md!<�Z$�q��0��q��I� �t�d�K}�9���b�ÛN��RfG)�����s/_X�2K��X��~�;�[�j�4X[b�^J�y�HN�ɔh]��#���ʜ���w7�>b��K�KU�T�*
��R5�?��`2eSZBS{�;���d���b�?��q��M�Ĩ�-$����� �Dcb}�8���$r������qj��w��'�5����W旑�Pa!�3T�*��X��d+9V����@ҟL�{)-(Gp,�(�E�dНd��;��.{j�n�#DA�,4�B����(V��<a�d�\�+��!
p�7V$M@vS������V^�?aQ��X�i����ʦ�z����p�BOu�����dq+�����&R��]���7I�5y~��'SDe�|�kz�z;�O�zPb �;���Ƞѵ�T��H�ǻ�zk�_��k���˪>�p��J��h~�sֱ���cӇ���+� �$Z�z,��@�*1�[���N&-�������m�.X~Os�6�?S����8�J[�^���Ĩm۳��yZ����F��?�K8
�E�>�h=)�m"i|p�nƹ�)uq�����tj�j�{Y���[��8�ƴ���3p6�*z�	
a�4��̀�������F�V1���E�@ݺr������lࠢRq웉�~��`��Ѯ�`vJM�����_�6I�湉�$DO��� Z��!Va�6X����G%#�9�ܸ-��'{����8�a�vw��z���Ty���Q��e�g�G����B����������i���8��]�'�@]�0�VP@ɦ���t�^����}�fF����ƢCd,����k��q�;�Џu�#SfX�
���|��s�^��[���8b��/|y���?�Y������]�G1"�5�5�?)�H�zDq����t���ٺ����TNq�^�t�G,�L�U7'��Bu���̜j�63�����<׈�V�UE��V��f�F{�B�Q��$�����.]����gI	�v���! �jZ��o[F��J¸��-���FJ~n��eR���v��4!q�ߟK4�eꚊT/*��!H^��gT�����C�����V|J�'K�AH�G����Ѱ��x��{��"���n�1�s�󜺯-|�H��@i2mɂMWJ�b,�J~�����On�-$6�nVW/�e'�66��R���з�kA0A��G�k,iʇ�DW��ʽ�`W���`��"�H��-M�	�)$��]�ǜ��C)$8�S����������Nk9t��Y0��n�� ["�S�七�vd׎Z�b�n7���ۺ�A�(��������^S��\�A�1��X�̗�*�F/�嵛��[)ن�:�ݵ�%����c��wA�#�bwa���b�f&� � ��Z톈��Љ��z����s1F{u���+5�P:瀢�dh�h�8Y��@F�)�l�Z��j�Cx.��3��o�n� -K�/�	�Ӗ��y��-�ߞ�m��G���L;��=~,A�]Ȼ?0���o:.�M'-\%�����Dk/�w]�=��RD=�bjt�l~;w���D���T& o����=�o��z[}���md
H7�������"�O!j�~�O�v�Ҏ��qi������p�V����M>�yo%s���ol���^=�@���~��C�|���7ZͿ�󥇽���t�-���j4�z��O�&Dƅ�R�y��b���s�.!���z��Z��u�!&��8�J�&ǀ^_�kH��C�1<���u�g,ADl���k��~��ᶷSD��Cm��c��ܬ��y}.F�
�`.�X�֪~��g�'�a<�L��2R��X$�Q�C��5D�dd{�A��\��t�N�E���\�;C�~��h����Y�=�4����]_:8v{E�Ts|�Wm�T��=X.a��F�®"F̛��߄?�!P�9F����iUI����h�{*�A��� ���~j�~tȜKC�,��#Ν�!����#��R��.�Cd*5����9&l�ͬ��ʄU���CW�?�������SZ��bv���.Ř�H���2p���,|<ZW娽���4����ɽ�3���c� ��/!���V��3�h��&C�Ho0��{���T�Ӄ��n��t�W2>����r˨ĝ��C��� H=G��~Dr�����zg˔�>�xCS�>�Oꑔ���(�mSȝ|x+��Af��l;�$/^�R�A��'ﲁv�Όj��6݊?���怘�Ge�7�?�k��ʕୋ���	(��"�'�D���$:���Mf�uje����5���(�\�dv�`��_1[.<�!�,��)Y��Y9B�����$����>D���>�Ŏ���TA�rZ���6�頾���L�Y�u�,�M�M�y<�Ώ�|�8�_!��i���I֫N�ظ�
���~�ړ����)湇!)r�Ap���ty0�n��:D���P�%]��~e[���C����wA��apg����L��y9�S�+_�E�0��_D'�`�:m�|�5���]���FtZ�������p$�d���U�@uf��뻲x2V��R�棥�y�8XY�`�.Z�K�Nt$��
<���]���<��*���������_ct!�W{��$=��p��2h�3ú�+ �"B�R�ly�sc�O(#���3>�i��ϡ>����f�u����q�&�*A1��ۈ�
�A:��.���߻R��i�}��â��\q�U�݈��8d�gQ���q��#T�j�1��77#�;%�����J��i8?U����B5��R�p�=ׂ��'�b"�d6��Vm�U�3<��TL�c�3Ƃl�gl)�b%c@��[��i��y�/����}������}-���s>I6;<Q�o$_B� ֙�z�0љ]��x�{�B6TǖM��ݮL��^l>���a�Ұ�\��1�ao�g�+c��� �̤в����l����d�̮�N���9M�lu�ko��Q�H������UF��E�t!�=5�����|C���d��tбRYno�����-a&�G:n����ڷU�ȼ�~;jj��(#k6�)41�ܷ7���hpx��ؾszT�����|Q�Ŀ�Fg��!lF����3 .��b\*�1ѣpw�Z`�3��tBU}8.7��\eY%9PLm�CK+���#�)4�}U&�$J��C�sa��ª/to`��TPw��꫓fp�GM�{}Bc*~�3g��n�OT�%o���)��C[��Q�5.J���mu�3@�=�D��s���y@�B��@p�{�*��V�}J��)nb��do��3]II���8�����9(I��X�:Y%���N��|�}}�׹��K�r���3���<�/)�����d�ʾ��ڱ��!L_] �[qfo� �*�(�rf,��C(aט1�t)��,�x����4+�n��t���y>��+��r4��dx��4��Minb�x�K�f!�.�L����=hxŮ�{�k1ED='{Y������9�n�084|`�0&/	�s�2Q0�ʛ� �5W*J|b���v�x�f��`�'l���I8�'�rn\��<�=�EB:��y��VRΈ�c�N`��i����pр�F:�:���g�-���"qr)���Y(<�R((��6i2P/��?�<����p�L�8{�9^��p8�sKj8�-�Do�q�l�������W�� ?����M�7S
h$j�A����0�X�!�U�>22���{�w�enP���o�&������i1��7*�{s	~j��&9���d�S9�x��~Հ�2X����$��P���7��}�`���W�v'�6cm��Sc>*�x�#�Eyڄ�5�q�6��ع3��O[1�]�� ���{�rrM�ޭ!�����﫝-�b��`j* o
�N
S�݉���-A���wX]�����ņ�N��G�a��g��J[k��@Zk����yˏ�6s����-�GY�3�(,������#��b{M"2����)܆�_)K���z����\S궹S"HTI�2,��̮f@�nH��xM��� �|�'nxϚ$� *�8Qr������%�����"wRf�鹑�j��k����Ͷ�T��������D�M��p(~0 �4��j�b��B�^���P`>6�̎��
3�-�,��ڪ2�y%耇��\�il����묮��̏��[�+�"Z���L;`
+�Jx��O �cѥ3���Bc�7`�V'\J���_���Du*7C�;��L�g�*Aa� )��퐢g��yЃ$�c}��o��6�2�G
�re"I��4#$�00;��P�e��9Y��cJ�������bsl��Ws�����8��h_���4��pLpǟ1�T�/)!;�I&,�B6��O%��Mf6�ʇDQF6��n96J�+�k�O��{i ����L���I���bF���V{�7��Ub)��>W�GHh�P��^{��C���v�_x��ah��X
�6�2��F���T>��]�-İ-�Iu�֚Ds�]�����k����dhdҭ*᳣��)[����Q�1��xZ� �v�������<B>�~�{��=TA>�1�ц�0j����� TV �B��\z�����^0Ldb��L�&�K�\]���;ӊ!��`��k�C�e�
 ��^=��v�����������w)Kb��?���iv�ls,F�#0P0L}!�#��=n���/v ���X�,�qEy�8?P?pf*2���$���?���� �s'u��JGQk�K,�Yͪ�<������ox��CL�2|1�ԛ"vb���p�	ʆ7�����&e	`X�����I*D(UM$
j����=`ֳ�+j���oo��*+��5����z �X\����F�<����5�Ϻ]x��uՆ �MУ1J-���0���{M��[.n�iN�0M������&����>μ��pc(q�{�&������M�n�F���xPZG��F�߬-[e�����"��׳�Qێ'd{��F�J�£�R,l��:c��C��g�.�;��E�-�s���"��)�[d�6����}5�Qkj�`ངM�r��!�l��Y�>(�tM�H����k<��(��Yt�'ñon��'���T�sc���3d��H��7����id3R9��o�:�֯����"ȕK	��ꫴ�Un���2��
�[#�if]=���:����h]M�b�<�x?Q��B�i�Ӳ5M��5'���J��v���s��,�c��R輬NPb�nY�M�9x�*�)��=E@|0bø"��>�� F�\����"(����v
���,�9ѸeoX��Xd��7�?�Oy
�<��Q<�8q�)g��!h�A)$�x��$���̗,�Ӝ�r�L�ԍw91�]G��{VN�Y��J��*��Z;��Xh�����!h�ܳ��6�\�#�tm���͝�c3�'
�&����e ��zX>��MD����]!߈�2��x�Y����}���z|h~^���ZTt1,c�\|�"��v��Q�e�7�B��"(�nHi��b�#�>�8����ةc�U�ûdF�vƔ�D���a��y�8�}d���8����uS�Am�C@)�a{|��K|D�%�P�]d0}�0�a��F3~��C~v��M�"�(��<,d�v��h�jB7��ض�h�>�s�k���餃&���[��T�H��k��lh�RKGN��k�צ�X��
-b��{v�k�HU_ґ��q����}k��((�pJy��N�V�)��}A�v'�QF~O��sfk'�n{O�??�k��h�C�1���]]π�"<�z�g1	xr\�
�z���Â�*�g&�aPf����2�Z��͂�����ʐַ8�7���b�����
�	I)��L��c>�<K6Q����yK���Y��C���>`��
%1����#�&0��6��y6��p��LF�^k0��R�p�#l�옋��j'7�G���A�N�r�������;�Jԧ�'�	�]c ��u3�ƴ_ *~>�.��ɖ+)����)0xdϱ�<�j�qک��`�Mբ#�5�O��D��?fFp���R���[7ҾJ+%m%C��wvs$z���{}&K)��"x�*ڻ��<T�4R�� �p���Ք�
�Ϫڊ�Z���r[��᪯[d�U�t���!u��Fo�������/����p���l�&�K����r�LL��1�4�.�ra~�e�|�yQz�\u�Զ��q6��פ�P��+��g��K
QP���W�����@�3%C�C�#����N]�|�J�#�	>���t�����iX��dk�:�w�[���U�_����y�{wfN����{G�|In�]���y��y�S�9�<�Gi�l�7��6���XI��ڦ�E/� )���׳��5ׂ�xn���WT�3̠����z���&*M(B�o�A���u�D=FwS��#[��*f��4E�R���zp���h'���+\qR���or�����;R4�=1��}��^g����ئf���7��Ŭޒ�ݟ�7O ǷL�>$�O���)�Wi�Ze�/���6�FΏ7�q�<��p�k:��ˡ����u���ZM�}[&c�[��A`{�� �=:����|]����Oy�U��r���Vs��*��hy�����x���L{Ѭ�b����j7AE�A�d[b�X���6r4��]oT�	"�R��V��_'��*��Q-b�U�+Fb50~��e%j�׊*��}���i׀@��Nm��,�Q�*[�\?�y���������n�!Z[��?oم	g"o���9 �籷��tVLIL�|7��b�:_p��P�<M���ڸ_��%m�A~^o�d&���R�=ut�sM`å��g��<���Z'q���Rò\3����	�������ng�K���FE��(��WW�ߋU�eQ�׫+�]���(T,���֞������ާ��3T�P�資���	�M���1�(؉uS(�PaQZ~Ey��慶a~�H'2[C�����nr#��b�iV�p�6�ɥ��h��@��s�|�B�aς��N��5+�o�X��>V��� t�H��oCiqU�6m�g�j
=䡝7|8� �˴�\3��Cq�&���z��=`8g_�`.Se49y���^�f���I&��C�
.�GLR�����:�I�YX����x�:fc�uVj(�\��L�[���
�U��.���][��)I	4=�U���d���؞��tpW�^���_ԯL���2��k�N6��t�vz���"�b�I���jn�ߪ>N�