��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�D�:��[괔�������o�.r�@ ¹�cr�{�T/bo>��/���m�qюn*k������WQ"����a��i��f*q}��od��ow��.8���0�8�[?�d�U�4u�}��~#���?<�
��VqN�jԱ���ـ��"-��.n��dmta�[���.�r��8i+�y2��e@�gC���c ;^y����ʣfY�E#	�j}�W����vu�0xNv�t�-�dV0����A3e�n(�$n��E	�
�W�^BM;��[Qy,^�>�M�ud�pO�%��^�lmFjiJw$e�?8et�oH2fV]�_L]}�j�n@e�j�?Θ�Y����J%����,30V�'f6���/.�{�!���ҳ&fmp���9�R/[I�f��ǘ{`1)���j��Gy���t�K�����t@���N}w���{,�V��;sL�����֤7����M)��19�x� ���܅���jh+���:����8B��ܿ���_V�*e�{^�"q4��t_���h;�{Q_Y屝;��:m#Ж|	$I
@���Ag �o����	3h��}��uX�&�U�+ٙ�B�gt-MdO�s`��dR�f��妘���}b���P+]��F��!�`0��1�-��^�D�Z�uG���z,L\y^�w�Q���4�����Q�惈SZ�gkb�17�.U"�?b�}�&z��c ���f����0�Up�&�"ïW�%j���Bf��	L�윅 �Z�q��	�~A6�#ۙK�x�D�@�7�%�n��@	F�����T��Em��4mx�J�ژ������Q���9�]/�k�΍)V���:/k� D�3���.���d8~�(|� ����,��c�s_��J�+����Л�旲���tГ�e�&əʎ��-��aŊ+���o�UVNL��3d|���K�����d3	��?��C��N����%FP��]�"�h_�g@9T��B�s�N�5�U�ﵓa�P�XE��f�,i��q�'!������,C��^r%���M�?�ta5�YS�D<�@���2����ԝ���	�(y� ������5��6�!���g��٤��g_��
*:(ݴ���ϊ4��M�X��cu�8�4Z�
`v��Q�sɹ����6U�:R2	0+�rq� R`=�z����q�
捒��� ~��@[�k!k�x������������3Z
D���4�����\V �C>�����+�yC@��#�%�Z�5J���=�,x�_����a��LK��P�"�j,P�c{q�eIo�6�x,}��1!jO�`B'�!�(�:í���������^�b&
��f��4�8�-|"�� n>5��Qx-�J�8 �H=�1g��:� ���F�Q/j��å�Z!����3L�`��>N��th�q�"*��u�+[���� A���1c׽�`���p_]�2�O��t�1T޻���z�B\A�u����(��d���A3-!	t���&�8V��v��D.��=��k��ѿ���5�e�Gy=B"�������O��5k/���G��1�
?5�-V������B̿ؑ!�q���L�6 ى��.ϙsT� �?�(�Q[L1%�����q.�1�pv�!1�V�S�N�l���,��k��f��c��5`�qS	[4�.�ҵ�ֵ8�-EZ������c��I�1T.��/� ��ڎY��h�)ql��ke!�|�t�ŋ��&
� #�h�Z��w�����3�^�a� 	��$���� ]u�˛�Ձ
�$��ĚF<!�s6=!�9��x�՝EF�|�bq��x8Zhn�G��+i�������"a�x��m��T):�ȴ.�78��Sx+=��$�+�6.x5�U0���S�5'��pS,��������0VY�D���y���3�����A�~ה�	"���Ak������J�|�C0�����g�J;�\ǩ��t�`Ս�~}�{B-<rͳ$�i@0=���ԝ+u�N5T��?� �~��l���֬��ن� e�>�,�{]�&A�4j�gr2N�{u�KCa�K��^!���l���K��w1�B$oO��t\AŔ'��ݒ8�t��#ZЫ���L�؊"K��+`,����Hf<-�a�= ���ܻ���o��=�8�H���_i
�tN[}�Q�	�u9B��n�)�춼����s���+��Os�
�[LaT���yG����Κ�>��L�?��W-��K0ۧ�^2���:7v�B���1.��
}r��=�*��"����bD:�VG$t�R��*�Z����|ђ����L����&�L�s��ɯl2 3~�*��Yi?G<4-1pK샣�+��d#j��Vi�˳n���g�ȅ����5Ӆ�-|$������]u�T+���K%$�y6fs���г�#u(�#b���<߂A�R���A��4�e�(���5sI�[��G��"P�� w*U��.h׬s��5����hzq�!į�S��{��� �����>g0Y�.�p���#���{9P�?�V�[�����*/��Y�^]�g��975Ǚ�\��lq���L�x�ˉ�H�8��j��
�0
�]l逸 ��gY*���wnt2����lBH�c��,Ỷ�غ-^~T��#�K��B� 릚L@������뉧�ʆ���IhS2�H��P^X즃ʟ@����������}B�%�-"I�E�����pǱ�8`X-\k%�+�Κ��N{|ڧu3ˣ_�$[
��a,�}���u�{9+I�ha�1m�yx�������ŨFw�������|��i��[Q�����v����������u����R�ש���͞;��7G�"o* �Z{R��� -�G����8��C�;����r�?N1.	јvH�	���
A]��A��'~����E`Jh��L������G���=��Y;���!]����S���C@�!�&�eNUÞ��c_S�����^��,�9-����aU���a�XM�j�D,��Ddd7-Ъ�=u��Gw�E�t�����Uj�vk�Q�=�e�x���ғk���Io�a�
+�d�	V�)Dp�r�Fp3a���}(�28Rv[�3V����)>$I �\0��$C��r�Q�n�<�=Qp$o��gB>�BV�HU� s%{�����"Ć����>;�7��%Yq����lHv�I�f;~����3�ut��k�����Wf�;���+>P�U	3p��W5J1/$.wu��s���L�i&�f��%�wj���5����I�8�(U�UN��.����>�7e8���O	���-j��h����l�w�/�~;L�k��4�(]��Y�v�H�� !��"Q�6�v���+rxn���c�YK��^3�kh�!	���+5&J���6���yM$V-���� �d�փ�WE����s��Y�P0���ta*uV��X�i�|Fr��^���u:�E�D����K��6{(V�oE��t�1瘭�b�G��,��kWd�"Bx?5*��2�h;�[tIt���<��a��_��y�Z��*�,:j�hR;N��؝��q>`��s�Zk�֢�)t	��z�k�҄|��yTYv
ɡU7ލh�U�I��_�5~nP��M�f!���T��DI�����}�&���U�#��퍲_�>�"������#eYQ�A̎-rl�Ǽf��V�pm�F΍������%sx  ��C.!?_��3Z��ϛ��b�D�u�!Y5,��$�Ј��R�L�+�Y����a2��E�.{�?X4�u0<����&x�7X�� �@��
�%��"r��?�Ao��b�%H���omO�����`�>���z�@�~�G�p`ď���H�oB����=gG~P�|�:t�r���V�.�"���DȊ28�U�Rr,��
,��ѳڋ,�Q�/.gi�9|�ږ{洍�Q�P�c!7-���@F�j3���'�����n�Q��+���O������}���Sq�i�K�􏍶�Ψԕ����tѮ�=qR|�\�-X��J�v�����*���P�>bq+�㸏��WqN��S"R=���/����|�i�x�� }#�/�;�+
▶�Ժ�Z�hS�*r��Lp���F{��2.K��!�<�Jy6�-�������Q������;�-\X)�}��e��F���߬��ŃaW�4�[z�ŗ����s���@���@�գ CDy��s
�s�İ��|�.��>�ͥZ��݃/����)i�?	��w��ɺw�"�E�4@�b�u��{S�����_.L���Й�E�`�
�����J�����'˥R.K���h�h�!N!����fz�T����|�	�?>;�����ɷ�_���Z'⢨D�܆vF�2D< ��7hN�~;P�ֻ�?�Y��<���c#�hk	vmB��җ;�Qa&���v�71��s�g���m0K�J��V9��L�>�(����XN��}�~ქ&K!��B�Ш�-k��@c.���i���?�H�^d"�((��ލ�ѤW�����NS���߭�)��z��F�~�?*��B���� c�h3��C�Z��͠���</��rM���x%�v�4�;�*�@�<����?|	+_L�sL!�ɜ��9Jܥ��I�
���&˵j�Un�[����C˄����@�PrR�u�����6(�-wl��)b/�����Uߵ8��:�Dh�>Z��_y��-�c>��C��gr'm��z=M�d�O$��������n&B�wRڰ�e��޹>���v�}/�B�'?����*�O�H�|��d��$��!��Й��:�����w��ni�`bVL�� )C���� ������!���~ɴ*������Qpr$*�"ħ�%�E+��] ��������#`ϱ9�]Q�0 ��3��	uұt2�`�I��je��*��3K*��AL�j��C�����东�GRc��B�A�V΄ӟ��'v���d����6�}<9��`�j�"���L���4��%i3j��f�ٙp�
�<�!V�*�3��4�f�zb��3�ę���)�jK��7�r��R��8�"�;@l~�U�uj9���6�5�X'Ý��\8)g�MPQ�����h�mD���z�j���Hre�~��)��bQ�C.��Uۘ��g�DNuNi�^`�p��z�I�X6[���9a4�{HD�ˏ�c,��x�*}�i���h��?�+k����ǋ���t��	��u#z�yjk�/����0\�v��6Ru�R�'��ȩ�xo�>L����sW�Q#ơ��Ϫ��ݟ7�of"�HI
�3II�����s��)�r݁(�caJ�U� �Đ��y!�	���SKn�d�(0`b@���A�E!{�$cgQ�m�F�(�8D�i��9Ö�%aQ�U��s�u$��N�0O+���+�c�P�24�U$�6�=���8ö́�T-�i���z�"{kG�m6��3�ڗ2�����Ѕ��� ��g���Fabtݢ��d�z��/��`5�Z��z4���%ğ��d�ߴtm��r���l���_5?�m�Pfl�hh]"����É=��"�:���g����F��Jf�Fʣ��>k�a�w햙9��S7��Z%\:���^*f���V-����U�ϑ�k���(�}��q��Cw��B6�
�A�_��ϒ��_�L��Z�v[�)�֧<��˧:�����9�g�:`di���'�q��k���{�9���X�w���f�1s�$����Y�$[��9���x�G!L��	�|^�]�ws��ed�0�����j���1�8]o�п�z���^��Z�A�1�c ����!a�ԕ[�Z�<�#X��X�����,Ǣ�����6X��z��)�HJ����"�n�M9�"i���Xd\33Elmb(�O��DA?)Nz)#�0��\�k����7��x��'~�I��R�u���=	^B(���{?���E�4��%|J��������e����~���(�Y={�C� ��T8�#�vތv�ۘ�=�a,�l9B��;x1���O���bbMNw��w����5*ZtS�(]ݥ	��&dǡ��!�"��a��.���ֱyU���_s�����h�<t��!�8F�'���M�}+%�����e;�¹�'(����ԨD|$(�{&���:
�/қ�j�[
	��(�%������9It�����X�>���<������`�<CVo��xA��rmN���j�F�7�\��M)Ǩ�N8Ŷ�5	A�Ccj�0��i5��
Ψ��}IpJ��DDW��C9�0�}��<c�=D~�$B"����?&������n�?_>I� t�U(#^���-��bD��sF��M�f��U�~2���,���w���fmN�	�H�����>�q؀���!e<s'>E��7��n%]��ǽ�ct;����=/�\]����V�Z���w��n�;�P�~�c��q>E���^�򤞶�ӹ� ����~��4�>����
�Z�oN'l8fh�Omԟ\�����-C��-V��盒^��P�g۝���XyC�������$i��`a��i��"uD<iB��5��g�$���\�o>Lc��7~��2�ڭx�N}�����O���E~oN^�?ϢZ6��#=��i���L|�w�)�z���;�!t>#<�+cg����?_����"�1�?sK�g����5�Z�f�^�*s�� Y|�����/8�{�
�?F��h��J"����x�dڵS�l�������2Ԃ@���լ�I ��ÍI� $��}��eLraB���Q6������O2�7j2j	"ƋBU�]��l��J㫒�����<��MH�����̊�Ӵ���P�����~m�|�np!���Rkl���7$\!�/�z��Η�b3������Sv+_J�l�$��R�3�]��n���][��Z���2Q�"0B4�!R��Wr����^��ީ%�O�H�w,Fk���'`dB�<3+wm�L[R2��],�����c��Cdt���lk�L��s>�a��v�;�@�oD�=tV� �/kx�&y�spo�Di�Y��8���D~�fn�B��ܖYala����?@锳'�41�K ����dK6l������a��G�ĥe��HN�QE�A��ۭg�Ԧ6�������E�0�s/�+!�.mZ9W�X�Jk��K+Г^���9���@����;�b�� ���8�C�ꬿ7�&	�#��cq�� ��q"n��9�\΀%��`�n���6~�"��h7 �^Q"�N<V��'+��g�hq*z��8���9O��7*8a��Y���{J��6B[-�G��-p�V�d̕d���G6�$m��H��[�42o�aB�6�Ȓ�{��lK57��}(VP��2�קW���-J�o�eC�R��a5�'4�}E)4_[�z�I���aI���W��X�H�&#`�c�R�V~g�G�/5�j���Wke����e��:0��$ʛ ��)�is�q�b]n�232��K�5b����)��IQ�o>r�Pjgm�j�Ϫ[�_�S$��� p��0��s�y�o���R1�S�!�K��ep<��^F�띊�Pv�"+��j�u	���j.�j��i�)��[�:	cߤ�!bj�M�חc?0�6^�rO���f_Q�z��f��'�K_�ّ�C^yk�R1;�u���P��x�R1�y�hm�����IC�ȝ�0�f9��� }�/�'�]�]o;)^C*�H9��ϰ��yX��Q=�bn����(;F�ޢ��,��4Iŷx�;�1�NY���,�I�H�V�%�˳��g!������tYO��v�6聞0*RW��2�
���{s�����vX�ϕ��绊�t��=V H_����72��\��o�Aѷ݉�z���E�����%��UB'����Kۍ�P�1���8~y�A�էW�͚��*s��B^1���SͶ�2�����|�A>C�U�H�L���|~@�����-J�`*wCD�8K�ϛ��B�^3�E_n�3&ۨDQ3�B�6�ݠ�{D���w�g�ט���{�b��l�OH��Xa�6!��@K?�֒"�0v����NIOF��O��9�[R�rں�r��t
��ѡ�����f���E��-�M�e`7漚;8�����b]F�o8��Q��Յ�C�x9��pp�b�x�R|��ב�Z��H"�[�V-��T3�vv�t705��A�O�=
�⅍:�
���n�
�i��ߙ���I(�a�B��	�L��������aiy��q��쭇�p�~<q&�;A����2�++�'^~�;Z�T��m�]��6�˾K����8o�5j� �1_5
3n�hN�3���Щ�H�b"����}U)�8���f��O��4XCCQ�C�HK{��dO����J�8�^/,�WA��J��%�n�@�P\׺����i��� �p�3�n�a�jV��<* ��;兀ށ��_�-`����[�_-	SB5�βi$�VN9�_�{}ʙ�K%E
����M�pX}�@FNH���Gt��>k�7(�~���tlf=J,�TqS��Xh��Z#���8bT���Bŝ=�4#������@j�Ju�e�v+�Qͼ۩��_z�2�A��E�b/���Y蟀y�X�9�O1��f�;��ʙ�]��Y!��i�=�P$ݚc�o
���nP��]�<t�0��o����bge?���рD��DJ��l(��X�ڲ�^b��Y�A0�YW�+����ܑ�>�0|���Z�g�GAL(�x3�(�`~?;`d�����]�L́�F��5�I�#	�Nz�[�|�R�T^�n|�:k���/�t���(�v �#���)\�q'�4��}
ts�7;�Uh� ^��H~�~�W�Y��
�V0��'x�\S�~UPR �b��X�#g]�$k�U�i@c�f�:��>�?ʦ�����>�����i0�M/C�.'�Դ�`m�ph#�����Ɉ��o��p	�;g���V��0�i�ay��|�&jAe���QTB�H�w��`����zbI�Ne�rY|o^I���}��m���&��/��ѭa����FI6`��/ٹ�.U�-���ڴG$�<��"��'JY�P3f>~ �,�H� h[��.FU�[�D���Ng���"{�?���_h�K9�_�`R8uT(�Qc@Q����l�Y��:�+9\+��y��_{�+?���ǔ��b��|Y*nP*�)�'�+��3^�6�� 6��rQ.�c*�e.��9DG���x���9�Z������n�rF���6�U6�}?��@Z�W�~���,a+�+����[G�j�3�|G����r�5��#{_�VF��3��Bj�%�e�B�˷�X��Wn��O�UƏ�r�ֻo�<=9�^&f�x��Y��N'��a�K�<�p�~��X�UP�!��zqz�sG�����'ߍ;GZ���)�Z&ݭ�`�	��'W��:@�#O��L�&��׺���^��	&"0�mZk�;�,G�5��j�� ����<�"3^Tt�^$ܞ`k��m�9�~�¿T�@�������zG�A����-`U��c���*�����,���.)��H����[R�_��wI�c{L�� �ϔb����p�~���&9^�$��[\Q&�X�Hy�Ĩ(���Bf�՞-q�e���h�� ߺ����K���g ����^[�͓���W�O���y=e+�"��I�[FA�ͩ� �%U�<��qxo;o1����tLj5s��o��y+��_�6�;?;�4����������[����K�M�i�~�xg��x�Q@}��n�{�v(�Q%�	��8��g ��	BlQ��)WݭBC�XE�p>/+�b��)d$�i�y����?W����"�5�gL:�7}7�1Ȧ�L��6_�Q=_���p_�(6Y�8V�.��}��@OjC<��E^��1�9��ݜ�V�~Y�a�`ؼѲg�b�ҷ�w�n��m ���M�P�dE�G=��\�c��Sŵ���Ȣ�&>�w��V�+�DQ9�����,)��<�'R��HB!������^���B�/�L �+�A���8���%�Jڎl:��b���FE�w���^u�!�ਇ7����+&oT-���j�a�!x���h�y9��ԏ EUa)��S�7�b�����O���9�Tg�"�xs4�$��n�"������v0C�_�v;Jm*{rG)%�尺��w��Av�6R�/*663��&j��K�}E���~�!��d��qG5�
�>�p}J�(>Y<S�؇�*v?O}�?�:��oI�u�m�tE�D��,��˞V��(��Uy�)U�J����$:�/�����1��R�K���:f=H��x6!�V	�v��.�ꡡ�;�'0^/G^�v�V�X_,���4�Y��Z����\0�SGp�2�����l �z���������N���Ų�l{�	`���Z6�?�W����0~�=�Q��) w7��8�j�[��M���y$+�[�^��Jd���6{[ʡ����K\(����c�a����9��Xy\�~������W�b�N �R�$��FU�)��w���c����A��� =^�W�x�7�}�������Y��Gg���Z-�j�6"}���
���I����-���y�L��C���Mԓ&�҂�eD!%GsJ����hqP���Vm�;M��>3�s��������k�I%��� l�n�;7����VK�o�J�$�\�ȕ�"J_~��4p 牚N��.D�ۂ���6���1��Cb�6�ʚ�xk��ɛ�������e� 7�K��H�ށ�ߜ:�W�͡Ȼ����;��Uq+s����Sƒ���R�%��m���5r�eL�&�!�JN4��O nuM��p���/�����؉u�L���xQ)bf#����B�n��'PU _MqVy��h*Z�B����O5f]�a�~�G�y�8�6�����46K[S�ao�vNx���M0��e��/i��ђ��(9�.ߗ������v5=���SZ��q����50�yu,���0�.�~�5_��G�� �h�m����y{��No�Ls�D�km
��^Ɗ��Fv��S�g��a����2o'�>?j�l�GO��wڣAS���mv��;�M�Y{c�S������;u?cD� ��G�"��E�*1I��ָ�4��F��o�1��|1֩ޱPk��5�1�>����nb��v�T��bϖ��o��݊3����)C�ß8;t�Qޮ�qc�R��B@c�����`Z���9-
:��qަl>�,��ϒ&��:�Y�ڳK��B�~q�-�t�ߊ2���G�
���26�?�����9&ПS$��x�Mݰ�d_pZ8@y�I�é4_�Åc�h9j��~Kv�#�y��;�| ��E�q�I������)��� ��ː8'p�D.d[^�������mm��FU^�m��älER�k�|�����'yss�XCL�k'K�/��M���gyp.dAΥ]��x �ǷA���̟�lK���ȒdIQ�!$�x��'Out�:Zg�aC@U��g�q�|k�Wf�>���]��E�x?�p͈+?�kP#%�U�����|�݄7�#���ư,X��h�uK��A#	�E�TM0A�0P/�B��ԁ�b#��3a���^'G�CD} K�qQ�
s-r�NB�-s��u��%Yh��;��>����>���]KD�gMx �������F~��T�b(��i���E|=���,�5�ź�;���R�V c�8h�q �ֵ��*q��z� [�R�,�;˝�H��U�˽[��P��7�l�z��@Njܾ��J����%ճ����UwS�H�����%hV�#3��Ú��V�H�;��y�C��gsY�9���Q�����,>1:�Կď��%�f��Ɩ2���=%��{�����Z]|h����X���e��X|0���^3wƟ���eJڻq` ^��n��~K� c��CD�r��;̡o�fׁ��|[=��Q��OO�����0���)�ж<��"m����!�ļ9K��1	#��<�{*ي�iy /���	��M�/��*���{��s�C�0�̰�b{h��sn��
%i��U�d7�>�1�EϢ�[�P*Z�z����		��@�BL=~%�ō��7'�X��� �%NӚ��g�q�s�q2T�x�_H+�Bm�LvBօ�zove[�Cތ��Ĭ�[) S1�z�dA�>����2��c���� z��d:hz��{�w���x� ��Z(��\J�/#^��,7���u&$𸺁���5Q����i�Np�m Ё��X:����Ũ���ͤr�{�ώLqI��3X�=Ũ�hJ$��!��//�RX�q�/�9c�m "�?���I~��U�㡊�=�׾����I��[5a<��Y�9H�r��A��I�0��~��B@tlG�/* ��U	�Ķ��֩f�Å'��_��}����jb�+����J��t`��~����2���-�X!'F(s�v�>g"�t#Md�y�ƺ�k�w�'�5?8�R�?&yA�k�A`���p$�A�R2
~��˭�^���g��t~9�C�C&A�Y��>���[M���E{ ~ŢI���q5[ � 1��d��I����rL{�-�&��S9�0�}�s�1�X���6�b�a���Z���j�e��w��5&�_;٘�S}UN�ݻ��'Յ:u��?,??�2,Z��C=(-�^�)�S;0,��$I���{.>�a�)����4��M�'�D,��Xɷ��Z��6{=͇'pp�`g#��| ���ϔ����U'_�UVV��H�{Ld�����r����{�m�	�A<]�K�O�	�.&Ł�N�G�����]0�	e���3��=��#*NU6�s��	��ulÅ��bh|)����4M��P��格<2~V̦�%g[�ڽfͦ/\W�x�I������J��Վ0ڝ�]{�T� Qh&�L�z�%V8���-��AK&�M�p���y;�᥾��l{3�P��Gה:��W�B�X����j;w{I���N3(���)ظ>����݂��S������k�0GK�1J������詵R�UT�W�I1f�<��m��Xg.��am�wȇ�UxfXZ~�1tI�����(�(��F�7��@�����h�Z�����Z ���$D�b?��{t�xROg�����,�[@ΕIjJ�����v�ۖh!AX�E�GR>'����@xd�τ*���ǖP�'�5 �f�Z㥳؇��n��/�\�r�wC]�-�00w6�y��꣜/j�M�C��G�k�E�ܲ���=fP��_�Y�=�؈e�u��g��Y��m�7t�6!���B��Q��U�3{��Z��3��/�M|��� ��V2ٹ�sO���D�pE���9��~x���Cs��*㰜�OCX�}<	
AӉ��T��R)ǛEޫV�G��'Q-�ʍ��7�10�=���Y;�KƦ�p9M6�m�ۦ����>�![.[�^��D���^^��ɏ�B����	S`d�}��qtK=���~�lc�iZ=b8�������ov�b�A
���"���)%}BT����B���z������;�M-us��T�[:#�\yм�ۨN�W�r��j�U�Y_j�n���2�V ��f>mGl2c�N�H<�q�n� ��WQ�yh$3��#ic��p�Q�ܹ��n[�L:���0X�G7]�Y�
�J!h-�I�	�G#p�����������͟���.�,��.k�H��I	xA��|�*-F�8��k�
�Xu
�f�t����.��R���:���;酭餞W�Uw���<�m�X���c��-j7�)��g��\���c�XQg8��̶���PJ|E+e 2�OȾo���-
.� �WK�fŷ+&8(�[�Y8o�2�"���BNr	��x��5���Aj��i�74#�%I� )K��z�����9��>
��{�2����ё�E��t���c�!�b��f*J�}�-��F/ũ��}jTڥ=�cO|�&Y d��8Xj������oږ4-��k�.�f&���	�^�� ����I���M��ojъ�]�)z�Ue��d|~�eI�~`i;R�է΢����*�fp�A0����u@�9�����b�tH���aT'�cr�� ��8QG0�%G�2-�B��Fz�qEm���w��!j�inT$�Ņ%y�Dc���A��D��UV�o�n�9	e/ %[�"�GqKU��҄EV`^��qV5��1n>��4	�f��x�P͘�1�~�Nc"\B�<���6.h9Q�� >�^��3����m��@�U�i��$URAњC&�Q�jM	��F�����
5���[��`[�6)c��N��V���>G�R��ek.��l��]/�ڴ�w�wt
lYK���$�Z;�̭���$��ʮ��2
>�@fȪM�o��#�Q�z�Nd}���sy����t%B��� ����9�\�<�i�<��lϐ�لU!+3^Ȁ0X*9�}2�HhS�E��Z,r8�7>��E9��L<M����?o\cE��W ,���HԻ��%�=}�b<��2��btD�}9��?1*FLg�Zx�3�m'Ư5:9��g�~bwx⩐����hl�������it������En-(�-1��v2Ђ�z�&�ڋ�D��5M��,h�l:��|Jr0�%!?L�۳�������)�^H�/�XJ�"�Yq1���7En�2��'\|��Ē�K�9�Ԗ8��'��gb�*�B���h��Ĥ�)�	:(���w��R �F_�p�2�d>L�:�ײN��Mg�P��9��},l�D�I 4~���?b�k}P�#|<I&ʼ%��"w`��BbDK3�8�n�R�d�v����6��;��E��|=J\�=C��^��]��`�9��dn=�l��cP�]�P!�dt(�g*�����N$�ȵ������p��y�e3㾹C��b�T�7�')��(/��?���Q.�F�3Ӫ�$M�"d��O+L�g%��*��15�_�7c3W�a_�j����z��~]hpG4�%�DT�Kp�I@�h�F8�F?wp�T0��)�Ȼ\\z���e�颾�*����-)��6�-�����F������!i+��Ƅ�SXs���<��aPr�'�J�IO.�?P�L�`Lĺ��M�g��\������_�7�uF��H��pi�hi�:I�6�X�+������`�e��2";�g!�Pd-����%έ|O��8b9�~+�t�˒6B��,(q��4r0嵿?�+A��Y�O�_��1�먜�/�<8�&J!0�AD��N$kY���I�ozrg�+�F��}+��Ů�?-s�%h��oU�b����Q-̈́#��*v��0Hj��U~�8G��sas���ws\g�:�[�Ѻ����C�K���	$g���BS����f+��ҏ?����v�w-3A�j�bo[邹a�m�NT�@��0�e��r`m6��ŰWg�z7-ݿ������7<�������j�SUza��ml��Y��REҬGb������H)ߴ}[�_Deۇ��ˉ2.�z�:P�.�;)u�CY� �Zj�GO�xX(О8�Hk'P�lI~�������Fp��`s���_Ə2>vk�F���~�Ԡ�\s��È�K���ޛ�f�q^볼uMP�U��^��61��Sa�����E�L�8�������o�a7G��UU���J ��n�/]�X����nkS��������x!���	R�*��(|��3P���Յ'��E�S���=��w����>nifM"��uJ�)�����VB
�$�-U��
~�J$����ϊLs�עn+礆
㌳�dԔ�|�b�&�����ueQ	�*L�(-���_ȓ����nt�Z�	���K�rI������e�"��G�6"P�,��l�1�zF�aﲲi�~��8���g�7���S�\�rr�!Ŗ�
���Z]������b2��CO�Vu��2P\t
��#�|w�9��|d8Tu��Ͱ���}oQ~���#��nE���U6�z�w-�Yǌ�G��;_����vh��I�
���Aw��fȈ�XRE�=�0g�-�\�X���vYq�7c�
9�Q�4�i������|��.7*�87-U�	�^�� Yû��U�?qۿ�͔ʾ���Wb�p`�Y�a����d֤4������DCI�Irߑ`�� 5�B�����8�DQ���d��nc@����S�ҧ!�B�md5_����3�l�cy�Yj[�'�xx'S�Y�S��n3��V_�2�"z�X�Ǹ+D
O��Ӛ��)/3n��[p�m��U���qyp�	�4'��zz��^y7�Bܐ�§�A� *��e�JC�Q(A~B��0'<J�͝1a5��v{l`nj�������¸%;�.�,d&)�C$5ז����Gq����Gފ�M-��04��D��&�m�7��^L`d+a.v��9�5F��ڛ���C[��z
K^@���L�҆�YD��c�zEI��Xg�-���l]Y���� ��=�a�bt�=��v�Vʰ M@�+�v�)�;s+�	'�_R�}��\�����=;#;1e��=P����ʺ�&��9IGL���<�4����U��Zg�.)�
�8G)'�Y�(�qn|�\c�Um�v#��
	=s����_�����0�����9�=�݊��
�:f�I�+�R8�-�O�k��?Df�%�Wk'@�T��W:�ۣ��m^���9r���
��_���x�L:2���a�OЈgn�N�� A�B��A\N�1�d�Sŏ�6n���W{�+�o�y?'�q�"$���
�!RF��y�j�A���F/&�A�l�7�L��8$�7�o�-ܳS�ּ�(��L�`׀re��FE��	�K ���pӲ0��_��*`���A,�8�uLS��q�ИD�ԋ*q�Z�y�L��+(���[�V͟xbr���5��Qޖ,U&a�ǍW���5^;���sV�Y0��V0�kK�1���Ca�i���Xk/ ��8�F�Z�g"����
�4�`��āKՆA1�]V����%�U�\�s:�a	�C#�� 7�F#����6z�o'����	gM���5m~�,�?;`�I��2m�n[��E�h��Ö��Y�<O��{�~��F���9vS�
6�eu�
&��Cd������}�Qs�߃����>�.] BB�52��ɫȒ2���f�j9��p��@n|Qf�e�����h�R|�"��z�f��܈���Ŧ1Dݿп�w��v[�����0���AUc�E�Dtok�b����5�'��z�v2ˢ�azYt�i����a�}wZ!����3���~�������������p��d��E����t�[_�3��g}��(�������I�A���X����?���!g�).ˆx��pJ�Z� S���0�F���O&C\?��+\�"BH>S�Ӹ��e�����<��Ȭ�ó%��Z�*_a��L�v���Z0��K�,��W�E�����E"���GS��o�Y�Y4�T�����	�����fx��ٚM"�а�d���o��HE�B���F���Z�Z���J뀕a���g9$Ķ��v���2#�<w6~r��!X����y��fG�;RuII�_
!���o��@l�7����`���-_�8�5|BRRL�����:5��{��4(��k*��&�}�0j��*���e1�Z�:�QU^��$Ja�H��J��J��71��A2��/,S\�LB�?/C�	���
�)Lx����q	����<ߞ2� �m�#��?�/��Q#.!ŀuL�>���ǥ�]�N��sR��~�x�+�F� Ny��Y��F��%x#ҧ&gh�7���'��:Ib�D�kB�S�u~�����x�-��%BH�{~�`4")�},҇� .�"x���ΌV<�
OEuG�ݪ2������_��M"���@�n���v�o��?ri����n:a��X�����λʬ�V-�.��O��o ���uq�T��b!�ՒI
�F��t��c2&��#�)�2G��8���(�D��3����3\+F����!חG����t�jy�4J�+�G�N���~S�ћ���
�v�e_�2��A*�Y�ǩA�R��֜V�����e��ў�`��=��U~��Wu�� �v������Ber~�EE�V�q�T�o����V��Մ�@)xl�k�h�~eqg����M~��(�*���y(DQ�t�d-^E��9��W)��S%��!�U����2�;����� ��XjYo�Ag9gTX@��v`��Z�|P���kϥ:u�'V�%���v�q�kE�m?ô7dQ�����
$7ۗ���q�ME��[�2M?2�H����"� �\����eV�|�%��`�����FC�W���~әzD�H|�=���}��Y�����&!�}��HR�P	��{�|����3�Cm���ًk灡�i�7,�
A�fs6�8c�����;�5�����@O�N=� ���籋�7���s�1�r���I�f�b�I�mW�"$�L�vx��s������xP����ջ�6߰�茸.|�0Z��b�7�񤼼�\Щ�?7ݱ��6��]M!����r�����6A��c\���(I�W��)+�� A��o����J�a�taN����0�r��x]K��ǅ���y�`)�����\U	��_Q�?�$n�q�hJo�N���8����5�XzL���b�Hu�Pu���.�'I�2eQϷ����|�hw`1&t�I�F,}t�#��'��K��'Ĕa7�����;ڴ#���@�-}�UKM}E�������*ĝ�Ћ�m��<��ȁ���B�L'`�^���5#��_�W��i�@
�*Ԋ�+�N���ނ��iR���\B��i����WuV��(��JZv�g��S���*�#��&p�Yb��	�lt����\��SC��K�Ǹ 4���Ņ�6R���t�6�� ��`8?�^sA�q����#����(�2�( �n��Y��q�5�s\��^ݳ��0�I��H�щ��o{�oċ��MПg]�N�*}w�	�����A�#o�d1�C�A{X�Y4DV�:E��-��U��O?�s�\ת�Zx?/,1U�o��H@ȟ���OF������3��|Ͳ';�	Q���>�e��wW�O�I,F@ ���GL/���r�����t5�bف�EB�s��r�b�U<ɞ2��
rӚ|��st�t