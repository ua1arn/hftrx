��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^�h��T���m�[�=�U8�@�|�}���//?�f5��[��M'a!�,L��ט%�͹%���K��PŽ���ߒ�����L�}t���f t<�l�h�Ķ0'56\�� l�1��6d���:�|Rb*����Lj�3v�yG�u����Tl��ɲ�e��G�ɉ-�=�\XHv��KZ��|�O{��G�р������W�zL�:����-&�H��ծ������1Y��RP���5ٟ5���<�$�zp�*1y���32	�;wN~��4�#�sy�+6��Ƥ�|��zѮ��lND��>&��x�s��I�5�׋I��qyz���S!L�հ���[�W&�R��hDPC������&���idowM?pb�DG�
rE{0#L��7#�^\/f�=4�,�����זoL�&vC�c���M���Ξ޶a.h	�b�$����U[scyg���u�x�Ӛ�������8�����I����P�\��H���!GyDB��׵B6[�Y���ߪ8q{��L9���J[��=g~��#�Pnq�,˗����jE�ɻ��V%Ϡ|���vo�/w�{O�ԤT~Wt>)fy �p��,��(P&�=�8�J���"o�� ��W"��E���(���4q(����e�y���@Y"�h�U�	"���[c2R��|�ް�cg����C%#�:z�0������� �[� ����^Γ��?�$<���Je�4���_�ܻ�.��`��ߒx��c(�?���B�]���;дx`4�|Ė�RVP��x.���Ad�T�D6���,kqʤ+A�bU�����'��������z��rS�N�����R5v�����D�ũ������g�O�jU��FQ�;�g����w�)��'i���	U��Ӯ������r���j��0���+~�e��W���vG�Sp���2�"JY��L�^<���O����Nr y��E�\:E\t�YUg0�k5�U�"��{X�%ĭKk�����^��y�_u���E?�	`6�*���;����Q�����iݢ���,M.��l�N	��Jk�i����}��t�^�F�R�&h��rrR]YE~BɅu}��$�;c}1h��
��,�K���+��s|��nj���o��b�.�}�s.�Qq2HP��"IRd��)Qќ/3 �����'�ӃC̬�yH���)������R�q�@�k�eҶ� ���>���{����
=j���U�υ6�2��u���>���f��׸$9�};H!v��\��BU�I����mF��#�_�<c��-�8�=V�b;�84��r5���Ƃ����6�H{�!��w�4�ܡ�.{X1������,���b��\�z^ڋ4_�d����������۪��G�0���k�d_�Bm\���'�P) .��m�9 ��6�xp��N=�ђ��U���6��]�k5�������s_^U�plX��\|�ۥ�-V�R��V��@��-W"��F���2�(�h��)��� ��+�d6��Lc���Q��QN���Ƽt�
����~�7���y2��c������j��h��!�cѐ��۷Vy_�/�����
��;�[7�iPj-M�2sy˙v��@�I J˺�!���v����.[���^�_
�۲�Sy�]������dRl����!~vJJʘ�5Q"�h��ӂ�;�V�fw8�aԏB1=@�i%�V�b�����Ya��D��sou�P[����44�I�*�2��Q�e���n!��G��g]����	b�"N�2��:��7�H3��2hu�X�g
Z�c������
�m��sO"�!��bFh���r��(��Ҍ��Œ���₄��bz��F. -�\�J+=ls!���������fd�\�m�p8dl���N���qؙ�ndIB���Ryv�'?>�}�jR��[#�n|^9pΧ�a2��ψ���{x�xf��"��濧�l����>��_ܚG6�<`��K�>��h�o�"0h���V�z8�:i�3�b���V��!�h�$����Њz�V�9�2�
��n0�� ����$+O��6A�����v&�M(�ZTr�f�y�l��I��f!ѩ3��{CĔ��ac$�ez-A�:��NV��ğ����T1FY83#��Bl����#��G�˓6���{�M���e���Q�b_#园�\�B{9 ��z����"���xP��l��������nqpf��I���C�9X ��u+2R�@h���,��۱�!�/
j�0u�2A��E����8`��Gd�p)��b�<�XZ=%߶�=����b$�3@��т�;?|��6����Mj�xWӘ/�j�0ˢ��=�28��@��j?��T�X}'��OaJ�N鐹{0�e��ώ����2� ��b�tC���G�Ie���cQ��d���Tk�a#���i��AߺYR��҆�Q��V�=oM��@_ţY�]�Q��ڥb�Q�KJ nJD��XP*i�rŗa��'������"����Q귎֓����ƖvW\^�Q�>�?������ϙ�	��H6W(m��{��+v���P:մ�x����~f%J��`j,�c��q�A�N��D����m�L Gȕ��,�l� �E����s�5A�(�W%�SP1,���}f7��"
���\,n���O����'�'pֿ�g�N^Ʉ� ,�p�I!�)�)�BQ�U�x���m�x?����if�[s��t���<�"�eç���^�٥-L���u�Y���<E���ʯ�ZUw�%�w�P��r��\Q!�W��O�wRF�H��j���Doh<�����C@;��NIv�I������߮�Š� `N�Y���������SH ��0�-Zo�oع��3ɷ%{��t�5���� `Kě�~o8[E������|�z\!��c-�]'�G+u���xE���$
��I�=�4�s"�D�t�1��Yz�BIx�t2���U%H3�?�Տ�!R��W6Գ*H侌2��Zz�~����M��?C
y_�*Rm��I]�x�O���`��r_��J�!����&���#����W����#�9����p�7o��K�o�*�ۙrOx5��;�gk?@��WM�4��=�&v
C�k�[f>��#5P��@��s{�O��˼�
N;HUs`�����-���iPĤR�H�XnǑ��Sc241¸o�r�{BL9�F����~�'�:��.U��Vo���w ����q���ܱ�4ܻ#/D��;
U\�%ӛo����U!�E5���.�B���(1�U?r�CM�'��=�D�6���=�Zbɧ�J���O�W��Z3t�$=��5q2{�g��-��&��F����,��2g�절hA��L���&�y<���l�L�`�l�bm���o�_�:]�}��u�`<���̾�Z��>��������_��n�,�T�(3Q���1��r�่vh�?P��(l�nD9Y��!���q�: ���e��|��@tk�)A�44֯���N���z</�м�ɇy�(ߥ����\���o����_b@�9��Ҏ����Q�=�G�ߐ"����IЍ/1�a ���c�u ���m�*C��*���εW|Q]�f@�,�Xd8b����gŎ֘���ݐ�����8��Q��y�����Z�\�ҿ�T3wS��3w,DĄ����f��`��̝ff�j�߬�o��x݈�[`��\{�UE�k�������%��nS��|��1�fNU%ƞL	�[,a�BM&�gα�U� r攩�6�5�F6�\�=�d�5@�K���l)2=�#�"Iy ��p���.,��k�	�	���ݼ�xQލ���w��t��²8>KOe,�R�`زu);�$�'��F+��M0]:#�!6�X�L��+���^�V+G��GFA�pqA�sU�'@��x!SfV%��0�zX�Sh_��y����� {�+_�C�(��@�dj�5'�N�'�!��S�M}7� �3����3��(]4c�:�� �<���8�r��+�z�����[��^~��}�;�3�;:�!�;��L8�r�~"}�V�PTuc�l�����y�j��u�%��~܊��Acx�	޼_�;�j���T�њ���8\���&��x�3)W�7"��.����~=SQobx�
��y��NiR^��&s��6�[,��屚.k�wO_;Xr�=���|ISߥ|[��LJ��L��i5Q;똋�m�.H���$o��*����E�������b�t}-�'���?ȅ�=w�\(p�@��5p��Y��k��<��1�sl�o��^ueJ����x�?8�c�E��pO�q�_���p<�֊Y��(�c@S��K;�{2B���^ڤ�Rg��g�GR�s`I�������b&�ּ�ȸ,����E;F�`|Y�1^�),)#��m(��3�aִ��L%2�����V���
lт�1{��B��}���z�ց!�rg:%�Е��z����� Ψ�$c��nݥ������)�ͫ���ŷ�c��;��(������釴�Y�(�i�|�5,2LZ5��Ϳ�����KJ��;zp���	w�Īdx���
>��J�:�5��X�������-�"f����+v��	��j���R �H����L���媵ͣ=O�4��3w��Q��"5�`<���3]/���aȔ��� W��x�)$�	�4Q���kL�5H��xY��O�e]�,��6�,q����&�Mws����Np��\J+ ^<Q���3l�X�rf����'t1�����-ܱ[��e���'%W�@~8U�1|��a�*+��t	!�&�9?/?1��ܶ[`��ͥ:�mR�ښo�Q�>Y,-z��P�/�$�*$��އ��~��L��1g�C��v���S���ʷ��UV]s��";��I���]QK�*��J�b��g�6�Kau�R|���J�VY�m�'��/�^�:���L P�7�>c�zL��p���	f�+��.V~���6e뻬�Ńʝ����P8Ё�h�L ;��W�|)�q��$���gz��h>9Z�f���v��q�
uz���Q�l&�{��Q~�`���<�)L��)�����$sU%�]��q�J��C���"'ӂ��6sS_��p�z�ݓ?��?�f�Z�st��mV<�}P�o�VN�P����� V�ΰ��PA���<��{M�j�&h��)�LdMLw9�?�*%t�J̇�:�k��1�߸�����8T�����yˡb�igy���%��jw��3¤~|�v��W";�i�e����(6լ�s&6"%���t$��mQE�+�S=�� � ���D%xB2m0�4xq�s9I\��*����;!���~h�gJk�͐���K�6�]����#��b����LYkn�Nc��w�Cn6k��}{��`���	X����פ����օiTӐ���'����>�O�<bO��8�2��y�`�L�Z��"O�I6K�r=bI��t��]�N�b�t��09)�A(�f�a�����َw�ܯ5P"x��uJ��7v`I��.�a#���/� �P�F~v�z�Q�|����&�k�"R���Ǒ`��k@�ȶ��7mj�s��/��_1`�02]�S-4K*�<��W��g���//d�Y"WLj;ϊ"�@�Na"��G�Td�C��;V�Q��j��]�����"��\�!���"��g��w�t�?����	��opU�ii��t����E1�%�Ά���f�H�K�Nn��$�dmtSڀ�i`F�&Gj�b��׶9�� ����Y��=LN��ʷ�B���F������<�Lw�)�_簽���g~=��'�m���>�E4�q�.>�YG�a���Я��d�9r�B��dF!@g��c
j�Xc��ھ�z��It��!D]��'|���8Cf�uom��������Yqт���хU-(�G=)%\, �p�O��ʭWh(At��L� ��E���:Z��ykz�J��h�]E�k+�GK:f�����m��������aG7�4����ȉ^�ف�T���Ņ����
Vi���V�ۅ$���+0�J"�C�L�)����͏w5�gH��P��۫�ns+��6\����uN�
�ְ̘b��E��sl�v�����&��z���G�t��g�[����\Q^�!�Ǘ ���D9��P��WRs>;,D]&�0������_;I�>�Џ���&��9*ĠC0�S&��v$�p�E� ��y^�i��64�)AȈd�)[�j,�՗J%���1����y�93R`d;�NY0�H�_�g%|���lE�`]��>RHHV5%sUNJ��dY7#��m�0�P��c��R���+D�_�ܩ#��M��u����!���jJ�C�AZ���%}��^�i�1p�+��~�����35~��|Jb��ϑ��Ƭ��A�kٿ��>sX��qX���c�L>�u<�	.��`
���K1����d�M0	�,�s��,���?M\C���H�4��w�h��Odrj����s$z!��X�}��c�4KkfQy�1Ac�ҫLU��I
�\�>{�,�g��g{��G��i�P�p�E$�V�|�;kI�n�!͡���|c�򧬼�/���
4��!�vL(r���$а��Ȩ�A I.�S�|�sS�8���]y��m@&�INO!�,�ܳ΋�m�՟�"�nfv_�!*z�'�n�,ފnE����WF��W�Q� ML����Il��Gʈ/�<���3Y�߲�z�B���l'7�zc'0xG��BN�}�Wa�ca;�yRW�_t���z&��(�,����@��&�9E�n�=����yUu�)�ސ,�k�s{n,r�����g��G˖$J}Ӗ�#��+�����h�Ģ��|��
qh��m��D�ݨ��N� ��SLzH:s��s����o�Q$l3�uJ��=N���iU� >�{��²���,�	d�E$ۦ�
,�,&n�Ꙟ���!;���Lq(Ȣ��f�n�T�W ����w����HݞE���^U%(r�V��w��ɬ��Ud�'�!�͆b�Ӕ�Y+��]X^��i�I}G����	��{p�^J�N��5��bR~���:�Ȼ`<� �������ޝ��x���PQ6�����D�5�����d�7���g�G�%B�L�i��b�|K��$��ttx�:��xt��iÙ��g6_���TC�Qw���U֝5٣"}�������f:�r����P����Q��bL��t�Z�z|�H�;`���=q�!OL٨�0̊p�ڐ�Zn�<8Ǻ�'��F��_m8�R���۾X�uˇC�bȉA �m�����Xr�����jS�~OU]D��)|��	��`i<�'�!���RǫR�{&���Q0@�5�*$�0Rl��B
��2UUG�/;�k2���:��=�Z��Ҽ1iOi�@�6S����|��q��~٧��lÞ����0
�6CƋ�G��h�c��a����Q���@����N(��/C�x��j�8�,z�W�.�*��i����-1H4�O޵,Mˮ��eȱ<��$H7����X�*",�����*c$zʅ��,�/ȯ�6�EwK��*�Ŗ65����S)�Y�0�.�u���cԼ�u'̲k7��F�	�g��4|v <Ϝa�d��5��:���o�O>�K����/�5��f�@	�0� |"}�9�~PgNl�(��	t���|nz���f���!贳Zu�0ٓV����z%�p��0�䀄{H�q��cI�B�����Hh��_��Y)Y	AH��ήS~�*#a��_�N��t��`�O���(8���%y�k�	V�CH�%��Kf�ƶ�IO���u!ӃO�&�ײ��݉k���u�Ŝ��\+��h&�g�v�A�e�"NȬ��(E��d*;�e�Ն�.E����H�U����Y�v��7TP?X����!�D�	y��8��C6^<g�C�ш�8@�z�ivG��WdV��[��jD
H���9n���Ǵ���)͏gb�$f��F��G�hKI�H~U�N����M��k,N�0�w�A�p$�N�h��"��XZ�G��*VK��O��!	$����w��د���޵��-T:Dg�p���C}��ߵ��!1�Ūc�ށH� T��9���ڣ>m枆���H�D#ɉd�f�N������!!�9"���OW�Y+�10V�ghd��/�ƛ�ᙦ��QC�b��Y�G#�X�I��e&L��L-���h�[�R��l�2m�(;�E��V�����-��j��=@�X�8�\"q���;Q�J~��3��r�W��~�[4����FfK��1��Ӌ��\֫P���.����J��i=��|�F��$n��g7l�;�т��F<�Y��W�
X�K4yz�ON�.��y@�	�~ᚭ4uR�9<�izDo]��Z�F���Wˠ�<�?�C���JUq�0Wkx.ϳ�lRA5o3Ta� �����a�>t�Rp�#+=��[�9^��7Z��K߿̢��S�p;9��!�}��X�����w��YL�S6D<}fR|
̲{��{����x�fC��q�0l4�tJ{feB����b�Y�8 d���O�9��&�cP
b&��˥뒇�-�,	M��w/�
�5,��wj��u�N�7�TW��+��@c������tz���~�:Z���3��ژ4���!�&���U���F\#���BY�x�A:4�LT��{��m�P�̟�0�ڜ�n��l�!u���R�|^(�X����%��m�.?����<����s�h靖50�y�J_�����ci�yղ��z�4���
���/�%�x�i]���l;xV`�����-�5'E�8�F�l�j9��v�|9��Y���U��Irr���I�8����^�:<�r�D������1��9D�9,&�t ^�L��5�HS�O�<�>͒aD흇�=c�y�:�����g�t���[�������s�H�nj�Z�H��)Ah�jX�A΢��d�~�C�U�؁P����]�>�y��;�� ������w��A�[���5-Ts&�W�w�����_TY��{�]6�.���?����D?Ȭ� Ų�Ƣ3n��gB�;d.@�o0#�98���6}7
�f]�I�ٓ �aγd��<�J}��J?����6�Q�?��B���D�V��������?�u嶯�\K��/^�3m+n�M�,l~�΃��{�1Iݽ�?����]bI�L�ʭ	��|��kҢX(Yc}���17O*���H�$�f�+�=�Ρ�TR5RN8ȩ�MN�;��2v!txޕ<�����	 �� �PS�J`�k�����vh���]��Vg��ӐV���7��_��0�T.���'�0m��+\g����*I� ������_bK`Ց��p�5Ruɋݬ����?)�'��z��0��W��ۏ��Jc�8nԛ��AjyO�mX�K@+o�	��ct!����_z��
,�FW���?�F`��nk�+�@	�⸄O�����y��I$�>��WlG��-`{Z,u.e֕L��&�����m;Bl����|3�h&��W#��s��Ek߄�Md��n�cX-͛��'���c�=����]Àe(�2W�	'�dF�琪��2ܪ��V��ǃ��Kg/_��g��l��0����	j���h�wx/��&���n����m�ʹ�R�
HW���Q�ER_�� Py8�$���g�/��5�8�(�[J�r�!�&�tX��O�Qݩ�hQ���T�8�-��(�+"�4m�t��������R{��D'�|�&�����(`�h��o���cD�_):=X�|��}{�9L?,��t|S�#�T�6_��.�A�,����|�(�s��}���2����Ⱥ4���l�B���Ib�Ļ���z�������*���]7����)�6�pˀOV���[a�U+�:[f��tn�C�*nuf_,=o�;���U$�Pz�vRN���Ů��F�ۯ�|>��}�yk�3Yg�T�yQ>�,��c9xq�7R����O��,���* �x��y��k���� ��<@�M�����K��(_���0L=.����B A��+	��`%A����Nd�K�^�rg5ٸ�_G�ߐ-x��V�L��yǷd�NJ�q��.a&��j��`^�wV���s�r��zN�G^��C]i��A��"*,^��'a!
�"���wK�~$�A�2����y�R��1d��J�$wE<�1	�@�s��E>�Gu%��06h)��T i��t7�(	H�/�/��l%v�G{X�W���@�2d���F���A�������UR�ox��bhrwx|�����{���%�<��>�����@���u��'��,���ЇlҬQ�'AvI�OԶ��M��D�V����V9\���/�0���#[��L��#(�ͦ���i�:���|�q6�sG�k;ZcX�v�Ѐ8��]_3�|�;�����	�YtT�me��%f����i��Y��W��$�d7bw������:y;�^O��wN�����^�־Ğ˟��a��A���X9������K��di���#�'l"#��f�,a8|eR�|:���w(����`M��O8�ׄ��o����ͱ��j�6�SL?��Ж<+2���-�&��'� H�˳��b*��-�f?�ylu��S�}B�W�ih?��G0�B.u@
9���?�l����Z��¾خ7���<&��p:�f$���]PV�,p/F)�O�F��AV�L�)�`���ёR�c���@�l[�!��X�	���ЀXn��؋���!E�C�#�)���Q��a�G�+�'nм�m�B�}x�β���kAr��'��l�-���~ԐJD�z `���/�������M�w�*�{&i��U��F<cG�-e>ot�a{�@[`�6���c���1pa�u:�ac��B.bO�M� ����e\��;iǾ����:p$���d5J�=Ȯ���wK����ӲS<iݴ����"�ؠS0G1���P��*)6��s�?��D	��Q0A�&�.΋�f�l�p��e/&jb�jP鹬2���3=�&	�ep��W�q��Mv���h�� �a��G�h�Nv�?������P8�	��b�!��A��y�7��
�f)�M�3Z$�Q����b̵��/(4ه#���~=��n�U�R����c�%پ���SxY/�(�D��0#�j��3zX�4�L$�]�ʺ��9E���ѳK����j�Zw�O����D�TO� �W���2�|��u���5-�<ᣒ�q#8�3�Q�t���-�IRȪ(�������.�7K�.��ay�p�@�j��E	?��?�Ȓ����1�6-�8S\�9�%a���QT�A��׺�B��F��+L��J9ԓ7&�B��%����a~ũ�
Š�D�P�gF~�޸KX��B	��3cz�kz�b~"�\�h��Y|E�&��i�MJ�'i�-����y�3���@��b�%�$ �Դ��}$�"-O��R�t#��~������&���-��,��;�^����d-6���^9t��Ģ`���xx��� ��ƙ�7'�q9B}�n���7g��~�L�}~��BtpV�GC�8���	��_��2+����������U����Ҟ���9Y�"°���+#��l��S�e�}Bc�K���!���aB�/�A�U���2��-����Pj��)����w�xGK��_��*��6 e��A_�����ck�݆YQ(4DI{b�����u�N~d���ܖ(��#�d�bL?�tC�_�7��4���v�����L�t�U���zJ�����`�ew�:GLb�!���05��X%��gyI!\���uZx~@&��]���9�Xg���3�t�o��u�c9O]�q�0��]����W�0Vd���G����w����/M��zrhDt��P4�V��E�z<Ȭ$6BY�42�.��¦]�Y��H1��B(2Z:�1�S�޺�O����՘�w�r��h�>��L��ōw�>����
U����lз�3uF���e�ݠ��S���鿰7�~����+{M�VbH�� �N��o"p7��N}m�{���_�oUv��Up�D������an����*]E� ��j"���{��H3�QM�mJ#0�ƲC��:�/2�9�F$�
nZ&�������W+(���]�5`����5X�{��_����I�,}���TU������7�=2� ��:�o��u�����2��̩r����4+_Nh�_q�Z	�IgF�0�{�{�dGgAD�&�M�J:s']�<�&d�B���B�!�b�N�&�8��V$��`�~�x�W��x{V��\���tk�SF'�0H%뺊Im�Wvv�]��5R<Q�Հ_R�}�5���{}(�"F���E�ߡ	xh;�p�A�o�����̮0��1��^p�|'�5�v|O�ٚ��3�E.˱^dﲟrb�^kj9��y�ז��i3+J�7k�Q�r(vە@���e{X=��� �J{���w�'DΌ���x��5�{�8P� q%���;��4��������VW �l��ӗD����y�+`��\HKZ��Xh�����C�U����0*O?<D�s�����<X�����pR�e��[U;Q���{wKR�p<ݗ΂y���H�������H2��y4~m���� ��{�6�f�W����fl�X��A���׎�v��`�X)		ĐA/��^�X�� E�x[�v#�5����Z	��?&&CH�x�Zn�ɡc�kU��`nj�,fE��^�ve;l� 5��51��A�ק��o8�F�5ģ�eȎ�ph;BĊ�	���P�����Ծ7%���E�I$!6�n�!S��~H%!L�z43e�hL�A�S�̿=���PڦSd蕶��ߔ%�EF�2ObZ� e&�CT��:�X�RXg�HE�Rh5�p�R%�ɠ�I���3O�K� �LY=��Z����t�p~s���,6���h���<�M�4���F3���/��G� ���Ww�k��8j#�g_TT{����%6Yjo�^��)aN9���9+���s�j?�=N�b,�夓�z��t(�z[�4H㚨���&������e�����)��.�[�|ü�I�\�d�;�H��}���L���J�с�+�C�P�g>�+�e�rd!���a�"z�p?vȮ��R��E{�8��z$y�KyJ��^�rُ>���ꠄ�nR�*F��=��]�l�(�צ��'�~���|gIK��Yʌţ�1~a�o�t!�,Q9��A�����W7U�1]W8���KW KS��o�8Q�o(����7�o�n��|!�FK.L&�!�n1�L/k ���,���L[Bx��N�%�o���~�����	�I�O�xgzDT�{��W��E�� ��ʹ3�w?���!٣v����k�bw
F��=dj��P����E�	ǵ���9�CCXM�Sk�҆���H ���<�4<�7q\�P��T��0,�)�aS'V��ՀXG�H	A(p����X��H1ɔ��+=��%��攣m��q6A��	R�߇
󵓘�/��ё� e4Ъ� �?#/I�f���נ7a%D����L%��И�`j��L�M0g�q\�f�	�p��oq��ӷK���ma������ax���}�O�0�\�z��ц���a^w�RK����Mx�4��y"��<�Rq")�^i�2f�0�� �d_5��bj��B�S\�����ը�J�~�rdpE�"8�+x�P����T]215����J07��an1�&R�f�n�Ne�rR�6��w<t;6
-R��`ܾ�T���q�>k�s��l�}Yy	���e�j�Z��/dm��j,�੏��
zdbA9-���ܺ���)~���C{�Z,�;%�y'&=2 ��n�h��j��"?�cdZ���f��\Ѻ���,3y��:�=4�����������W��qp�Ϻ"�U;��v�L�B�TI�}�~���5����\�a��r��^&��O�^^�/e��D�@�Au��e*��dġVΤ<6 ̸COʭ�x����y���sF��E�%݊����of��_os{��>n�����q-ʃ��[x���&�>Lp��\[�K57M�M[��{��BG�����9Ac����m/f{��g����#��Y�¶深Mf��28-v,�y)>{�*���N���a0��gG����Z!2B�?E:�ב	��;ȱ/������AI�;O��0(���l{2�_W��)�'�׭�A����аd��F;I[V�5wm[�2y�5mmO��E��_�?{��
�2�,��TW2my�B���6��������� ���:rR�ܖ���p�{�n���N�j��	�u/����Dp�K��� �;�R9W'u���A&3�2lȲO�ُRB�0
�6�=�~��ދQ,O����:�s'��ޘDF%��o���^l�����e)��_ɀ�����%����֌�u9����Y��%)<�]��ھ4J���o@[Z%-�P�Ac���]=M� ���l�#b�������m�����qW��,��hK���,�ʤ���D�]����#�������.�sj�m�6�\y�(�!�A��?'�<���(����x3���M�L���<���/����}���J�w�a�xR�3U76H���D����ϣ��<��}u�tZ���<�m����+�mh"Ô�q�S(�n�%�UX��vTOVRDu-*�F��"ME�E�y��(}�;��X�}��L�?l�#ӿ.�1ʊ��_��Έ�P���P��T�����W�
B�:��l2����[F5��hQ�V?��}m�0�P���z����������tن.J���tH��s�W�*
^+ɣ~��+j��T$ ��uVx$*{߷P��հ,HY���8�\�Y�"̅������\�M���P�?���ef�qb�/_��f��
u�0��"���KG?�"VB�k���q<�5Ǌ�Oms]�+hV��y)��)���(`.m/iŦ�$�#�WQ�;x`9��
s�!ɴC�/���f��K�x�`�*GDb�K���p���T-l|	�5�i��c�2[�Vk�N����:Z:vD"��M�<@��� AN�i�Kru���O�]�a���<;�bs�}�H���}�p���^+G"]w�s<3 �si��*��`�����xwy�Uo��X-�K��%t��1��	�q�+L��4�T�>����_�Г����;X<5��G5BM��ܑ�]�����7߼K݃`��m�^&Fo�����G���OMt㉕O6dR��L���ʒ�7��My��Q�N�A��QB�K���\g��/~�;�
_�>�_�I�8�$������*D68Č�<���e
��_n��@�R����:!�� �3�V8y=�ӛ������:&�D�%����.�9�3cT:9����|�v ���6O4�\�C�8�]��br�f)ktX3�â�%z��Q{E����Ew�F� �}��g9l�%j��?��@�#jB��la�tXW�G���P�u���2��\��+������z�7};�-ga�\u2�S(�Y�<�V���d���C���pt�yC�,�Ŋ�ќf����ʳ��te.�0&�=>7O���I�6�.d�X#�1ةp��s���<�4�u!�涃��s�۪��'O �O�塆��G��pL�
�[O*gR(����u��{�����a�ݏ���Ϊj�{��+�q:�s�(�ڳ|�SO��z>��19����SW(�r��?#Mx7��v*8HaE#��ݱ�����l�$��Lg�	��l�2D9�"��Qqdz��ۈFo�6��#�:���E��[��>m���������ZE;y�f28l�Z���n�����/4��TRuFg���(�1�{�>��K���xo(m���<��{��UN5Hb�F툽ю��~���G�j��g5sjc}#���+���Ğ RXH7v�m�Y���?$����Vj�f0��`�8D�(^'�_�}��<ê�]�0�5i�n��
�ljQ���o,��W�� u�8*�km��F:e���]DZ~��	>�	p#!�M~SA�I!�u�0D���i���W��)�Vc�jGHO.�uIg���u:�Zl���1�`�,�Q!n��(�t\!.)f�o��N�a[���2�P�6�H+�M��S�=p{�Χp����"�-!ɬ�T�N�E�X�����䉿�-i�I�ϰ�b�W�^�v����ˎG���U~mЉ-}���~�N;!�'��Ԋ�ۃ�C}:i�"$KKk	xͻ��-1�h��FX����Շ�^VS 
*9�ӫ����AlG+a3vZ����xiߛ���i��)�x��-���v� d���sK��:�'�F�J6,!�G"��֢�n ���%���rs�Fh���-�=0>9,,&��'��2�I�e����u{4K7C�f:%޺7����h���BK�hV{�Iy��W�d	b%4�
�Qٱ��h9B4�	���\Vyw��]go��Nf��<�mxdcmAt�C�����f���`&&!R?
߸�.⏇�M&Sfk[��n���U����j���1w�u����߅����@Zط������P�ED=����M�L�b�EP����� ��4T�b_���a���\� �Ê�p���j�e!p����4ȳ@2�	4X{A˪<��!y�ucj��D�,z�� '���lds���^�jOfS�GIK~Z��}�D���� e;bu�W,(R.��N�1�d)$o�blfb�B����4�υ��#xA�B�	>Cnl��6e�i!~�C�^��H�D�;14UT�bWz���ybq>ۣs�ED^���#�[���6;��Y�6����;���<vW��u�����мZ]I�o��lv�Q�9ʣ��Χ�Ftr�_�6տ�3� ��;Mr��s�2f9/��Z^L���k�`ى�F�s�l2�@J��BCǹ���|���k��5s���R}~���O"�"V���9]x���^J�K�	â��]�1��O���	J�)Es�dR!��g��ʲ�U(�P�5�����ȑ{=���̖���Q+oX⯰�G�S!��;�5�^r��J�ҕ�-�6]46B�-Y]3Q�f�����?�-/m�Q89���.�3�r����@~ɡ�.$]i�@�#FP��ͽZ*sާ(��@Q���'��J�����bpI
"�&R�;�X+�@6Z
|c���O@�IϦ��tv#Kų�2�%�j�p���#գg�a�p�ձ:�	4-/C����x����X��!/�<).��*�S6�1c����Hn[!$h�-2����l���=V#��YlŲ�}uh^V�R󡼖II�S��:���흭�k���(��-�Y�/&|�f��U�1K��D0fѼ����F�8���3N�bqB�t4�nz^�z�|��@]���Z��F�,���t�7`�%�˴B��Q��zݤ'��v�'�Aɠ�/�3#l=nKa��s��?旑��澩{h����aNvP���KjG�;И��������_t+O�[x�nqرh&r��{m���?�WS�G��#�h�X  �1L��0P��w~�wA��m�TgWa���eM�h;~���7o�6��XQ�e��D+܋��+���=}|�����2S⽌dW��NH��D�$�z�2JΡ�6�*Q�♼�a�� ��E1!� ��O�g/�
�)���g���ݲBy�!�|3���i� ]~�ɭYlJZ��������P��3�t�E=��ü`$_�i��o<���� ��(=U��_�hj�.�a?�Q�r�?P�_�,�볩Q� ��sU�zN�~5�?2vjU?[��y����a�R�PvJgY��i�E>��-�Sp+���*�I	�4��	��.���x����A˙��%"�+)���  e%��a�0���0��������mk":����'�*�\
����=�4a��bv��0yߢ?��`�L+�׫��y�n���9NK�LY���{�7��]���c��Rq���z"x����|B��L@'Ӿ�<�E��7�lj���iI�����MF:C��ρ�ޠ�m �7/wz���T�<�S���Iڗ}�����ޙ�'���[�!�!qt������J������b5, q��I�4-��Vv ����0U!���pX���_��W|�V��A1S4U��i���#۬���nJ��:ʛ��lg(�5�a�xA)��]3n[�3kU�%��(=���wK�JKI�z��b�v��	�`̲�i�Iӫ��>(�!R���$��V��~2Y^r?����ĈQl�]	@�=�:�k� +���-a	4a�D�IF��"ܹ�ߑ��7���F�����G�FY�g��Uv�!��G
o���9�of���[��	�lFv�U.c�ӧ�H&��)Y:��GU�
f��C_�\��5@^�����̤�l
�g䰱����ZHˮ�/��L l!��	�T.�t\��[H<%`�l�[�C�X��a�gd_[���'뙱Ry�Б$X	�'+��n.�'�S�٠U�q�O�������q����J��`��"�=!�\�Na��
�. ��χ����19�rԶ�Q%���w<iT^Ԉ���ۛQ=~���Q.��[��8��%��v�DblS:U�D�F��Z1{7*y�VC͜�(�gY���1&L��+�3^��v�s	p��#����aл���-��0�lvb�k��MySɊ�Y��+��K���ݔ��B��Gt�SA���%�E����K�B�[b�c`�A7~��M�>��9��7~�D�O��/�	t��E����\�����w\$�)&�SD�1qu[Ȁt�S0g0=EL���]�r����=A[����]) W��{ $�(�.Ao?�1ڃ�\������A�P염12��(D�c����ýx	�^�R1y�nl�ʱ�S ��� ���waD!q�ͣ2�J�V��V�����Գ=��U�)QN�Λ��ZR���QP�;���y!8��/��\Tz�%����:�j��L�ӏD��ua�t$�*�wX(E�w5�����@���)�u<����q�r暈�����}|�T�PB-6�"�;��s����o�.���
xr�cAlý�����-mx� =��%�>[?�S�*V�p�C�y�7�V��s(i>UG�+����<M�*2��2�TZ'���[M�ě�襯���rEAD�~�J�5`�/7�!����R�+��e�� M�W�:|X��k�<�zWz&�\�>ssC��%�4����iP�7X��ЖPX�ZL�h^wB�X0��(���k�tV��
ܩ�MՅ�$��eK.J��}p�c�Nl��VA��~9�aHI�٤�d��q�d����qK�w�C�$��Б��m��If��8c0�ڹ�gS;�8߸�R6�#0`���b�Y���#e@.@�5%8��A����Ⱦ�8�S����"�#��j9gO�Q}Z��M޴�r<�()ޡ�-���6�8�&�][�K��h�V$5�_��p�҉����&�E����)�_"���Q����^�Å~A���u�\�!eӵ�f�D�д�HBv�)������o�����	` $җ�R�o�=˫v%��'�c>M�;��}���M�ʝ����	���#ʊ�hr)#���ܰ��z�E���վIi���V�$�~s/ft撶,%����j}�������T��uN�����=&�+��ɹ4t����۬��)���c��)k`,��3^�?6��D}�bƟl>&f��tIZ���v:�w�o�`��[��壧Gl�&�(H�ğv���"n����9�x�kN�Nq���m���L\���*����"=ҷO�yG@�e�y�)�Cpo�~�A�3� ��*�H;�V�
�?m�B+T�s�BrNZ*�L�xY��Ы��$�:c0��s�Dٗ�M��o@k�p��u��6�������������N�������;�%�˦9YJ7Э�ч�«ɡP��a9��+/:���&o �b��Ȓ��@ςv�10�v_j?f[A����n�s*�3�r�o�ޅ:�E�#�������er��Xz�|M�vӶ� ���Ͳ?iL�_��b�1x(g��{�Z2�3ZJ �lyk�/,حs��S�t+e��1�!�%K�
�zm0�V��^��$�ީe��A�q���yu�H7���������O�č5}�(�$�AI����h?,
�|	��rp������i��ȇ�ru����!�!�4�C^I*>��6�~���gv��,��0���LPxt��L��f�s�8+���J̘Ω>1Ӑ\aD*L�bj"����u�R3{��>c�B�y۟��&d�N�Xf�S�=%,��(S̗A>��B����.b���j����MV�/����IߟԲ����!�w�Rxj}!�stU��,�4(c��tfg���qj��M� ����ތ?#ԁ��5GM��-�@-=�X'6\��"Fq��y�W�J���i)C&ce.��mC�@$٪!����N'���O֏���E��d�ո�H��hv/qATh��4��xCHq1Ef���m�8E.��~/�	�⦫Y�7 %H:�����
-�D��g�a��/�Z3"�����9�'�!����z_-�ӡc�ֹi��"+����C���oϔ����	^̐��u�o��A^�B	�6~_��%w�g�~[��]U�M�
eb$���%��ѧd*�O@1����`��V{w��P%�:џ^3���(�7ڳц��ѷ7#d�>�D�@��`�<�gع}ˍh��áHA�+�w�*�C�i��	;���I'A%t��ډ�"n���(�:0n^���
�sM4�C�I�^�,5G�d?h��X��<���?.�#<$$s5���a�?TD��e[?��b�w�IF�L�����9���u�U#�A+p ����(ԚeNN;�@��&�r�*�\$��zE̌�I���wC����ro�o����w��͍�!/�ͺ�'����`�Ȭ�ưl��C;Ꮵ}�Z�=��\�7�kp��*N7�,�j����n9Y�Է���|����w^5�Τ��-��d��(Y)Y*���V(1����;���-n�][;��ͺq��&����\��;H��A�K&�1�����H�܆SQ�_�-Ɗ�Q�p��d,}g��O��~n�xq��0C��s2���t�"/�FU��[�#U���#���������=�-W�N �i!	�����ӆ?�xމ�JZe��f�#��u+�ݠ����l̅
�Kp+�>�-��t �h�'�e�����[��i��1W���h[.Ss2 "|�ㆩ�$��5��z��c��qRot���b��(7�5S�� ����M�Ϥ"Z�u��p&[�}&I9�Z��>��#,%�h�n}�=�l�@0�i�YZ�ԇr�NߝcS�G(�q�p�H���f�* cáM�1�2I���?��������M2y4��VX��3��81k^����d�w�(�m���l<�n�_�����F�j�J���d�%���6���3�6�D�<C�y�"��`>VM���?p�3�ģd���7�H����O}'���hj�����Qog�X������r�w�Mgm~盈�%O�o�Q��&_-��� �x���G|v
߬�����>�ݞ�թ��\�|X�ஷҨ��%4	f*yz�I!��a@����ȝ�V���%����"�Y��x���!��������.��a��0E`ʆ+�'���gG4J��b0��Õ@� z����M��Q�ΙH��d�dt%$UU��ff����6L�������B]����?��6J�vj]f1����'�����`204�X'�E�\:�G�,��\dW�W�xG�i\Nl2��ܟ��*���^>��������D�MňAE��s���q����S'Z8}U�%ۃv���L�&�噱�f9ߑ�Gr��&@�C���Y]�ͷ��j(��YwI@�G������fl���4{�E�ݦ�}��Uw`�ƃ�eE�v�y�>�ւ@�M�Q���T{i���Z!�Ba	�צ���&Y9LUVw1�~)��A�2�ڤ�=��9���\(��}���,ӡLq����HgS��oe'�|8 i>�;��~��&���`���.�]�v�8>BϲJRv�#�aя�7���,*gc�qh�f�O�K�M;s�˅rn�<V¬�[V��iV�`pS_��y��v'H|�
�M�h+o�sc-LjwȮ�(���H�8��mF!�Ś�Λ&��]�=�ܢ���������5%��i;ۣ��J	��>�Y��2����0{=�X�[t��@N�WR�Ѩ��m?�R}o�`k"��q����/����0n[�kw�C�،�?�<�2�6�U�SĉY����C���XJ��>�p��xH`����Y��S~J�c��1��*�:���IIBm�� �V�_e�s��$����%�e98���ˢB��"�IxK���)��tf�7)[�-^x�sD w�"�<M����s�Yç4Ⱦ�7�j��������-��唳�Ɉ�9����6[��M�"O�5��{����Ũ��`#9d3��TԄA-#����鰿��:�s��foPJp`�	'A/�W��]iX��Acp�Ϫ�l���B[�^-��O�D�����Z�+E{9A�������O�u)J�C���J����1�{wM2�{�h�YB����p��zͭԢS܋�D��(+��䪈���ۤ6���!���k�¬>�1��,t�T}%n��o4]VM�~|,vd]9㻾��㴳��k�:�"���MZ!3E�BMzrK�%E�D�6R�{z^�P�(�����	|�o��I��~����_�Exܭ�>p�nD�P��J�E����Q�7�>~��T�*8Ƅ�T�87�X�s�������?i�x�	g"���$��37J��s�`i(�[s-;	�g@$섥��|&4
�d�; ��v&� ��:��&���$	���ç5��}�~-r=?W�GIٛ*���LU���Rϝy��[�d��a�� ���l2�c*�<V��=���B�g��|!�V����y�4��h�����G�?єpN#p��Z�4fs3�Gb��ך�� �8D<�Fl�����ʀ	d�T,���	j�1�s4��q�d�n���;l�޷�`Xt�iF����-?"���)�S��5��Wmsx �H�dn���������9m�&П-y<��1��u���>�X�mh3���2��X ����(.����b��wξ�������O�nd���V���`�x�G;��΃�;���vkX�/�x�Z�U���8�T#p)pDj�;��d��/:���[�k	�h�=]-�k1ck�U�p�k[juP�+���/�������C2���U�,�KN��Bk�Μd������Y��>�3D�*�����d%1�����|�JQ�MI��:E��z����ó�_l�S��ކ�L)�ƿ#�2�#ab31p��~5���F ̋����2��>�����pA���v�d�ʚ��(�T32�8h�AkU�� �N�ѝV}aK0*�B����H�s�}��)�f��;�y�a����_}l�Y܉���x��ث0�:y�8n�H�p3R��6��S������-�M���XI�.PHr@T@Ew̆:Zu\�b�_�jrk�ad �͵���q��We*T�F���O7fy0�\��N�o�͒Bմ�{�U*����W*���pS&|�rS2���nIk�z��+2��ի)Ɲ���X�`���~���SQ'2͙AĴ(��ҝ���u-���ɜ"0Z�@ W�S��X5�3�N����O�b�Pi�X{��r�Y2���i�a �%&+@JQ���zs��z���(f����Om�؇��qk�y��|T�B�&����S� ��jkrs�\�E�~�]�}��F�čрl�k�\���7�o餐w���xb�Z�6!��6|�Q��l�M�g3��t��K��j.�ǳ���'�튡����1������ �4\��cm+adn��j��mq�~�l��`�g��T&�./.ی7, ��68~m7`��ń>Ƥ�~HB�snv�hU�����Ɉs��������8�(u��\�T���)�n���'p��2�h�b ����)�Z�)]0���~8�$�C�>4��l|%��/� ����͉�B��S/��&=c7��~������쿎G=(�	��ְf�L��4>S'/��P�?�xcp������VϽ:'V��$�N\���8�!/V�C"�d���=<���

G|��p�sH�ʶ��B},V�+,��ODUGO}.$��J,%]�=´�vB��%�cqYd���	���MJ�ǃy�����C�M�S� LQ�0F����Q�e�P	�GFb��~;�hg�Y�Z���r��US`�s5ƅuW�=�^�N����@F�/Sa�f[�~�6��qg�4[�]v��z�_k�-ƃ�����H�ߓ�1
���T ��<� ȥ%7YŇ�=xM�7����  V`ǩ��w� 0�M%@N�AU�!e�Z@�o�}��Gܝ`�ɢ>�{�gr�yt����+���1j���e>�J�[���͗�����:3�<.������XN�G�ju<_�"��$Wj�@E�9=�s����9��;?W�J���~���,E(�b��ݱ�L�����]P�֨���{�|Ǹy�RKɒ���	�\�*�o5����֦�h�S:*��KTɒ�bdv근�CÙ#��K,z��&�B{_%�w1A��ގD?�j�v�Yn�j���t��Tz�TUᥧRa$���4���?������H�l����d�L$L��k��;��VhA8=�� �',�=��Cn�MO�jby�PO�� �)[��Kħ`��(5�fx"GR��E~�)�C�E��%�,���d�V�}�sMF��Z~#�,�Z��l'���%�4�I��=s�Ԍ��8}�Ul�zA �VB����̋RN>qj�z�^c`݇#+����1j�C9�F���b��W��ݜ�o���F<îr��6���Xb���CKy�C�H�"��٥���v�'eQ��qc�lኽ��g�9q�ɮja���Qbv��1�vР{0$�?���g�t$���B�j�$T�C񱒏Ū���?a_"*�	Lܟ#f��U�zm�@�?k���YK�v��1����{S~��J�3"A��ϥ��t�5wk�I��}#M�+�M.�$I�$�ML��?A�P.�� ��f�	��1���c��%¾Yw]�����j�*P�2��1��>�*-��HsJ�TX�s��<#�$�ޜ��W:=�ǹ�>q�z�i��Q���!&�C�6��^�[�˞����~w�Y��~>tWg���Q	�*��ck�5�o��q<��1Lf��b��@�j�`q
�s�g/�$��s��+���ۇ�a��� ��yrE�1k?�J�����;�F=��|��~����$�����P���2Y��S$�V�Ա[
>x��Ԧ"�Z#��������$�e	AJ�ʆ�T��p��\�
ʌi}�0ĕo`��*A�ݟ��s3��6����|F�|5�X�zwl_����i�dы}�b4�q�ƹ������a�����#�ߔ:W�58h3`�Hg�֑��K���Z�
������mɾ��3����?`j���s�=�:��WO�]TĊ��NreĶ�'[�`�c�����k���%��\��|�Z��D�ש`����Ȅ��#�0W6��M�
!$����{�<4�����0��T'>.g�ӈ;P�	�9�S�\N ��Ӟ�� Ws��ٝ�:�'6۲�k���[jv��0�K�!�V��S�j/��$�Ԭ$EN�u��k�K��#���JL�<��(�:ą�X��l�Ú�מ�<��w�u��40��|��p7�n:y�xs���K���I4t`Ґ9U:nq�#�A��Z��"+R�F0�ݦ� �4�R0�_,���d��0ߎ�b�>�uV^{3ڡ�C/�O��?xF$�r4�m�J��1���X)�
�$�|ȇt0�F%@����j�J��0�@M�RØ��������dn�(��OZS�L���ß��Kj�D�	� Y� �Հ�_q� p	B`y��@V�������;�Y�k�D4�V7D�.��s4�>����>�Ǝ�ჰ�Cn��\YUi�bU���r+������ه�>�����G������z�쌋ጯ����<�Ip��o �օ2�z8r�7Jd$XQ��=7��V<�?��̿�� ������F�*F���ߋ+���\�^��VW.���ia犏��6���JZ\Q�	�a�^�<S�YP�Z�$Z��}�Q!��Cz�Ԉ���ӥ��7�
�Y�3#y�ꉀ�6�z�?���6��ʉIm�,��m�������j���{Z*���4����q˖���F]���{{G����璘c�,���8HQ2hc�;Oi̤0���2	��8���'G.c;���`Ky����
0f���Q�7%�P�@���_�g��l	nաn���/2s��޴�G�@�=2Bh�oĲ텟����eb�ŗ�tk`
�	��D�<��z�XI�����ъ�|nw���0d��v.��D�ݻ bU0�(a�jZ'i�z�Ɠ<4��bo*���⟒�@���#z�A���]W�,��u/9� m��)��h���v�(�|A�W��/���R9������6�7�0Q�ׄ�����Q����ByƪC3��
�u�k���`;���Oȭ~��������Qo�K�*D�5�8P8��Uigl�0��]K?�V쁢!�ǐɭ9W���2�HI��ꎁ[ǲ(��+�(����0���I��q�^��L�MU��ɥG��j�£hZ���n"𖋏NBp�'�7��&�R��I�o���*��,8��s�w�P�E���5�ӿT����L�8��N	�y���HMs�T^����z��\�����!�	�����;�o�����C�}(�H��ޔ_� �I�,��+P�[U���'�o�x��<�p���F�q��Z������H+5p��U�mCjUǓ��]��8��R�~~��B�壼O\%�$\sBC>�KA�?����w3��8�0�l�Z�e��)�h5�z�
NB�}�x'`_�]�mMT�~��M �Р�3����*ƻ7��~�׳8�V\\;,Q)�oMb�U�Y���&ʵw=�J�5��L��8�2�6�Y��)�Q@g�ڴ�d9�r4
Zݰ����>�o����΢�`;/�~	s����B-�g�{6	�gʯL9��<oދ�~r�
h������mJ��^��u����P-֖~���E/m.,����8���o7�ZXƭ޻��ά(n�1;L,�aJ%�x��/�������dѲx�Q�v�||���h�Q���i�$ۿ�Af�N�nzz�8@�@L�(!�@���5@���O���1���� �<UC/;2��[C֥��"���=�G�2�Ծ��H�Օ;�2|ր������DȌR�;�[�F̥)���h�Y���Ә.�W��e�^����޶�q�,�{�C�@(0�t(d��ˀ�� %C��.�*���\_+i�Z��4jq�=���"&R�/J�`�,�H��K��$^H�W�������@6����B�&#�r�%gkO�'8�@�� .��䜃?�c�9�fG*c�#R
��<dARA�y�G���$�Y7o��x,q'��G)�XP����,�s�ӭ8^c�"M��QϽ�>�۩
�h"��4G��W��F@�[�E�:}�/bk�P�!�'XՊG��(W
��h$?IA���k�պv%�C��N�&�is���A��3>�e5�R�s�Λ�}0t���[���V��vϣ_���v��~�K#�h��Tϋ�>x���t3PV�]�� ����̑w��,v� �L��1V\�v���B���f@.�.�3�Wb$D��F۰[��sa�f�@R�7���O������Ϻ�%���Y�U̡&�7!v����mM�/q��#+
��|q ����P�kz7}��6�Ӛ=fN泦��?[4�V!���5�t�<P�WN땪����	��Ú5�j݁p/���h� !�2_TU����
c�rW
(�L�7�`�Bd�n�A�~o+���k�`��� :����'cW|h%���4U��(��7��w���P����
�'��-����UR��݂����yEr�,
��\����±^3�̩�_��@AH�
ؕ��`zKL�*_���̲��:�lYhԓǋF'j����e��]���@����Q�ZBs���4>3�B�����tm��1�F�V��R�B2��{��q�w	-Gm�A��{�EЗer(�ۭ%1��wmc�*��/�q{s�Bv�p��f��]>���z=qe;��A�L��{�@3zz\�Z��W�/X]�#�=�ۖ�r��vh�!��^O���f�	��t}�A=�}����2���D���*��QS^���!���f�2�,JE�d}1��Uݏ�Ҿ�\<~�˙���d6M�M�L�`r�zL�������=q����`�W�����%ͼ� 8@!��y�5l�[6�o��V�t|d̉�t��yO������@/�h�Z|H>�i7[B�G���O��0@^7��++8�G1���> �9al_l��%�?}��Kd,�������Zs�c��_y�7��^	"�S9~�)6�p«��W�����u�v�4�b�QJ����Cz��	G��'�]�mP�7>'����m�ݝ���Ŵ<P�IآM��6`�����A��`Ό�Oʹ��ٷ������JhNZ����*�y����z�� �����Z��ͭp�<
Ӵ��bM�F�D��\�$�<E2�m�{��iR?��%A�"pv"ȗ�n�]���v-ڠ�S��u3�ҫY|~/Y��W�+8�Z1|�1p�����@f�E��~4����`�X?�����F�R� *����ξ
��R̕������%�^�#F�0}N�'>��&�\ekN�+~�������W!��k��t����/���<���:F�m�)��˷0ڭac��l���=�Gyt;g�L�?B٣�l�׍�H�~����
��&�_��#�;��}��{�Y�ѥu��r��ږ�+F���-11��b���C�4J�+k�a�aMT,���{+�޿����'��}��֥�6ɂēC�󊍃{N�~�ʕ���[���Q#t]8�X�̨Q}Y�d��1�b���}Ҏ?P6�!tȫ��b����v���b�/�$t�\f^vs��gd����$��?�#p�&�8W�����q���������DQ6�%�쯘��[	y{��v��Gg}� \������Y�t�)3R�T���ٟ*!R�5�_��o�=#e����q����梍��&W~2n�bN,8�_�e�:p��.s����, ��eC��ݥH_�y�@��`���
0����8��F>��\�턬)���&�5S�s	2֘v�+����~�ڄg'�H옄L�����ځ�}bv�:H��Z�5�$8J<�HҺE�B֍�ǌ/^�s�h�k�z|�Y��ܸW��&�n��&a����Q�M�{I�R	��:��f��\4.�bٟ�eg�bk����.�$/�@V����0?�C�Z�R��\vQ�Y�d�Ih��{���PԈ)�M�2�#�dV�!n�ʣ�L�[�'�7.�S�e�M�7��k�y�,?`9����l�vf���D���s.YU���y�dE���_����"�e�QВf���q?��BJk ˀ�ڶt�n��)TVe�r��f6����5��<j��eˎl�iE �jg�J?"CS�۩�=v�Q��9wm�i��H�&/b~�:.����w���(���r�a3s_XS��AyM�q�!0
\��O�~O�;V7��0�M�8���vx��.���n��W�>���5��=�FZ���'�.^5^�^�:ا�Uhz�60�]���R'=ȴ�v�t�Nk�Ale�dx�as
`w{)G&��µ/G�[�abS�`�h�%�y �c����Y�_�_��O�_�qcT}�iT�44v�$kM�&� �]�f���\H�e��Me�R�8�?n�=r�'̥����!JW�9ߚ���k�G��$�T,~�<���F��9���y���2�kP� Ӭ����󌨖�)���|��� �D�\{����W�	�I`�����-yW̴[�(m�x���B#'� ���{�¸}�I�ih�y�j����1���s�	��@���&Ў
D�E#w��V�5I$ -�P���$��W�����	b\�lY�0��0��R`?8��gA�!�X�`��O�s���$�����py��2�n��|��d�x�}-�N'K9Df~��14T�8�Q�O�Wmm�� �����/���~-���D�*X�z��#GO�s�J����iU���;�D��\�}�����	ʱ���s��.���ź!kDZ� �i9��~��_�C6ϗ
�);��QΙ��T���*�_�~#��8e�e��/T`��̩�)�����|\��Cs�aF,�oh9��^���P`R�͙4hI̲�(n�����߿%���w[�*/�K:?h���f2��pX̯�F���I�J���:��1ԩ1�ss[�ei��N]�c�!�W7ke���L�%{+�X�l���.�sEz�	t����)��F�<P�/���{c��^�ˣq���<bo�{��o�.��
[q|CA��⺍|j�L��}B�t�����yM�j����wXt}6GZO����H_��+b��#�iI7�.�<�����^��N�&������*5�m9�ֺ��䅨�:wu�"X�<6q��� e��z2�$�9���,���|��ۥ�:�0O�.���O�I�7�f�l�ӕ欛zm���� n���O;ĝ��~��pD�=7υ+�i}Τ��r�[$o=����##\q9�p�R�r<���S�#��Ejo�[q3d9krF���w���˺ ���h��ض�S���i2����K�Pk��9�I���Љʣ�L�/�>��_CU�˝o���iB@��|�0n�T�k{�L����F^l�JƫYC���).aYK[��P@���Kb�'l�b�C������������ZR�;ʿDXat�����$
��9�ʑ	�j!����HȒ�>:�8�Y-Zw�1�f�����D^"C�/��>X��(��p�m{cre��F�JȦY!ǟ���4mпB�J��ǲ�()\�n��&S�U-���t�SΓ�t���{�N��Z
��FA�;G��v�(t��ƈb�U9��є����>�oT��<�0�llo���f<V��A�Ԯ���T�v.a~GA���YR��	�q�ل��S�<�@���><���䡴߯�a�dL�����Wg6�95;cج�0a�Q[A��&RT�����W�v�z�����V{
n,J���*��\��u�m��4�W�~ㇴ[{F(�]|�C'H)��u�47�PF��ХQJ�k���������i�����׷�O�jq}Eҳ��h�v���֭t�# ֻ�%Ӊ7�1�d@)������dQ�U�<�uT��.����~� ��w<�u!���CI��!�u��9FzFCl0�(���
��<M�py�o$O�����MD�����7�U�'S|z��yh]R�my.�5���-Bо$R����� 6 ��_�Vc��f��#Ŏ�1����tw|�~w.֪ RB����$o
@��4�L�K���ú�������XCCpb��Z����<Mם���N�����ri����"�,���ǖk�U#��1^z�:۔�q #�^���Su�+H`d��CTc�BN�V	(sR�cVi9p'T#{���;E<�/���~.��o�+s�0O'���L.1�۰����/����+^����lU�,���O9��Q�.ϟ˸����0*M�h�U/�Ú�}�t�R'����<��� �ǈ�Z�"�ߙ�������yb����|+#%`|AC�g�H�Hmv��ȳG��!��R��wjY��J��.,�od�%���8�)]msط֧�����uK:�x�Bx*�;��o+�~[�C�|�
y.f`�e:WȽ	���J�Fh����|��w�m�
�A��=�!b�3d�����<�	�������Oqpbi�8��B[�Wi��'(Fę�^?�����4�8�8����<V�_At簭��o�Z}���
�G�r�d�)�T���ݛ'D�p�-���-W�ս���N|(F�F}�YW��|_��n�0/q7�V&�!���f��r�v������f� 	#!$��-C6���{t>Y���v=����D�e�mtfJ鄐���h.Zيy>�b(��y��Iߛ�(���I���%�$D�+��,��;���Md郭b:��q���}$u�R#�#hܔArm!8=������@��,}��'�{_�X��*bf3�Ҕ�&M}��(�:��6�� ��e]H\R���������9�X�cRu�h�pP�&E�\ץ��
�ܔ�ӟ��Sy�!,����v��p3��y<_�M!Y��~�!?��}<��X�|ư���S�F��W��~��Ij`Ɔy)|Z�%�����jy�������E�X����Ql]�^��N'�m-��4W���v'���g�|/���5���gp֎�%�?{��{M�`\f&u<��g�YeKP���B�u{>��Ȏ�H*���ɶ�r�z da�8��|�W.��L��lx��}�����X��B{vmc- #����e�dIM'��u
����A���/'��U�;�2�;W������&������5���&�'r㫦�c�6�m�}x�;P�m�1����1�oQO&HX�P7x�2(@Zc�6̕�ƿ���uf�< �$�WP�e>?`ϑ�hѠ�\�ݗ�~D�&��Lwq����*�S��iwS�G��W4v�t�V�X�2t�j���U7y��q���e��;�(��xd��L�g�-�&�v��b�+����S�RC9��
���_�{���j�(<�wO���7����$921֖�1�ɑ����M�.WZ���ܷ��?��ۈ������B�\���=�>�%�E�}z��ҭf���q��o$/��g�P4���ဟ�iC�4�&����6E�����P�q��7�{=d�?��`��q�OD-�����f��o�y�N̆-�ଅJ{K�
�ې97MJ��8Z߈�%W�w}ҧ����+�1�ސɁ��	P���2���T�K���U2(�~���1S�j�҈�2�����eo%��'r?/rSlx��U����s��A�!on���UG���x^h��:Y�M����j�>�S��ׯ�OC[x�8][pֻgc�<D�f�5AI0�=�PZ�dA�ী�ޠ����(j�����j<�L�x�2<�?|��_�r�kF��	3�@���Px�k���]z8i:v�Fp90N�\�Р��Bڇ-vض
<�<��I���X��*8S���o{�;��1fv�b�
:r��3��˯o���a��:��_��XJ4{9k@�ѯ]��q�j�SG��m�ho�;�x����V�� �ˊ�M珫����ׅg�K>��� Q}��p�v���Q�OF4�K���8n )��S۾ؼ>���~�V{��6��D_�<�\� �$������/7�ԅNS]�po0����M��Jv���	mR IF�[}��0�iH+��� @J�R�]�V���DT�T�KQ�ԡ����d�X&�����D,��(h��� ΂`e=,k��=dAܯ��ʯ,0Bu>��|�ң���7�B�������kU����0�V�����K�#1����v�����\������4=����@=��G��䬳KRG0h�w��B�HY���J��X~&��X�a��1k$�~�k��C]��4t���A�o�ixжD��X�Z!��I��+�� ����1�ӭDF[��-��_F"�9�cU��q��PE|�JuS�'���}5��p!�ɥk�M��m�җ���a��� �fͮ�~ZO��"�碞�$["s�z�z��9k�͌#�����hgb_���D��R ���c�z!�e��#��؄۞�D�rt�#%{qH�	0TN="�#��È9z�&ď�'�E7ב�����Т�9��+T��j�K�XQ3*$?&7n�`���QJ�HsC|�xX�B��@��~�6�Xy�\]}��{ö^���kٺ�s/��i�,�"g�Y�+V!��tRP��u��(�`�5�?Ҝ�W��@_9��'�!b��]�_�.6u �3?��5�x��	��e�5aǷ�(��H#3���J���|B��(�)��2=�2 �A3���7ɐح��1�,^���J��PNq���Mt��2K���b�T�L>8�M���H*�zt5L}P��#��v�������+�X�z��S�3��}�ŵA�CCp�(�$9��F��7���<{����q�z1���XT�?��	�+>�h�H] �l�A��k-j�b~�>�'b��r��B�%�����-�faj��t5�v2��w���B���bw���]���4�� �qF���q�\t������&�UǼ����p���4P~��6��h"��Z�w�`�"^#��a�B1�����l��7��HciԹ�gA���&�-W��ڍ��,v6U�/����e�9F�Th�S����'����MĄj�('���n�X�a����S��sD��C�d���1�L��!���#WhK~U��.��n����|�/�R�I��Bl�BHabop%B�B�|�'<T��ɝt�<5�I��g��+̠��ksH�m�_e���d���� ����"�$ۘ��Ȱ�ȅjt���ga�jn)��&	\y�#��������	l:A��Ӌ$��i��~�p���{_��(�1�Z{ -�|pݺ�+R�)��R_�y��?]��(� t`:=�����Wu����]�nfA��R��6�N2:�E�$I$�٣c~�
Y�!��g��G�ep��٤HRo��~ S���fݔ&D�[c_%*|~BSW��8�kM����D�D�%����e�dGB8���c���X��J���}������ti�]_�����������(���4�t�So`�&X�M�/ɋ��GA�b`��$Q�PL�>��:x�u���ۢ�=���F��B��B�}�̣eJ��k.�&h�]S��+e�KMB�1�2��	&��(J~��B�ΞY؋�Ω��^���͉�`i���eY����K���6n��4��d���Й�d�z=�y@�ʷ�;<HM+7��34 ���
M� L�[�����^�)Z�74�uTo�i$~�h�P���a"��4��̒3C�.�
`�
��F�*���5��z�q&�����;�r�a�2��0�2��ڦ�xݙ��̸��'oҔkw|��4��.V�T�|�����&����}U��D`G$
F�!Bs����,���B����3!�u~O�vd�[#�k7� zA� �2+�|���6�� �o��O4��)w��,+>�RiS2ʲ�9�l8���AcO����4�����V�3L{��;�j����BW�C�����Kx�)�T�1��kV
й��
m%�\;yK�x8�$���&G?G��b���~94�g_e��^C�J�F�#1T�ß�u���p�kLj�u,���l����@z�\c���Me��Ɔ%u�Co
�眂��~�#�嘄Ʃ���V�i���9�{L������3��	��,��� B�}�֚hЊc��0Ƀ�xٟZ;g�B�I��^8h��v�s;Їl��&�Ð��U��ڿ�CJ���'�	l�$��7f�iw�(h��)�{�h.�еz-ۨ�TɱIܘ����-��t��I~���6aȵ?��:,i��g�:���[�v����rěFB���Â2+N��4@�T�&;�̐/ӱ`��R�����`4�.>y�m���M�����م����f�T˴<�n��0���JQ#d�@��
'�����?��R	1��x���4(���T�#�Yd���%!�̒�aÃ}ǎcPfp�������Q�����77=����|R7w�M ��S+�P'R)��n~W�Cx
��,|��8B��
�{��ם�iv������V��F`��g�Rm���ac��}.�4���c�R;�&Ι�K�$�����Q��,�9�bK��ex����˽�.�jU���{,>]
���]�J��F١���Xk� O[7�y�W�r;�9�d�aޟp,$�M��J�%���e�^�+��:�z��0��
����#o���$��}��S>�G� �/��D�=���~:'x�B6�7��38�pO�H�����'a�Kh<x��[�M񁣕��m+,�&� d�(����7}�KW��q���1�Ѧ����+���6����p�M�3a���J5�tfE1�d�l.h�=����C����
V�]#D^�C��'C���5�q�P��%�-���'��>�f.Pb]�Dy��heƄa�!�9�q;�%�U��'�	~p�~�B���Ԓc*��p'�~٪�H��bqQe�c���5"H�P�/PV�f�����I���X�,A~��	���|y�ٶsFϕ�ob>���$z�l�J�2��ܰ����l�2�#;�Q̌wi�iZVF�T�9���.}�=F��a�z�5�M D�{* �*��ˈ��Us;7�;�8IT���Wk(G®zǉFs����K4aWǞc{*�['�%��4σR�C���y�b��0ؤ�\��Nޜ��'�KQ�x�����n8�����{���m�{�6&'�K���A�[:Vb��`Aj�z�QEH��i{d�����ʑ^�~2!�;�'H&�J����٬~u�"|C|���٭��I�Q���Y��5Q�7��W�.��LРG�3��K�z��!a܎����:#$4�0�w���� �!r�.�u���v|NX��C������6O�i�G����>`�^:�U����=�&y�'2�ȤC��M)`����]�m�B�-~�#�c*�16:S�q��L'r3m�aM{6[��}(�fe��Q2�#$O�â��O$�Y�8`tw�G�çx�DC[/��r�X���\ޑ���k�{�ݒ���و��17Z�o}k��Ǒ�P���3Z𬢟e��b��}<���(З�+W�}
\�f|)�o Y�.},餜�yusl1�S��ނl�"O�ä^f7؏�$;����ⴴ���d�Q����ͥv&x�.�{A��}-&�j�QKpz"�xS�:2jH���񶩼w�#��Av "Y-y��9|��ҝ�Z������6���	�/A��̍Xf�t��,@���x{T��	y�cx��hh��O�u�ɡ'�+����h���U0
7BPf�<��&�V�"+��,9"\��� �[*��W����eی"Љ����a��G��"�̎�\A����JI��-[c��1�e���X�c�&C�^��̊��f��5�ӞoԒ�Pl�q�;�/] bR2�"?�h)>N4���ӝ���,s@=,��]�W�00;�⇠1a
��TKCt�����1*,����I󨂾��}O� ��0+��p���$\0���5s��y��A�z�GS6�[[Gg��0ʞu��"ݶ�aɊ�Ro/$`c?W�F0�/acmB��zq4���^wS�f�~!L�n�[xN�T� �^�T�M;m$��Z,�`�|X@+Zp:�~�~�C���s�{�]O�y����[Z5H���N|��H��9�|��E�t�x�q~4M�Ɣr"���D!�z^r�F�F��5/kſ`*��L�=����L��9��9MM�ɺzGQ���f������e�X8�	>�	���0Y��`*�~���*��Q�.�er�;�O�QAw�c���1B^�M�'����;��-�}9����;@b!��'��sV]SJ8��`�����z�t�P�x1q�X��	�
�b��_���{)kl�q>#�l���@����y����2��T�M�o��+�"����j����E��A4V�㐏Pi���W�E޸mD���R�ZƗ)$�Xs7Cs���d�G=&�wT�H(l�R�������#Q�LQ'R.��j�i|�`��$��|�v~�%����\08aC�k��_�%�!h�"}�bvg~��%�33�����-q闘V���ܑ�M7iS%F-�.G'��������n��&�ꕲ� �L,C{������%l���f�g��Fv����d�=��Q.
�C�m@�%�#���isj�R��)�|���UBʴ�/�(상h���@"�t1��o�?|q^5�T��9�6:�G�
uT*t6n��c�B����UA�OT�������
��Vy�+����w��9�YX:��x��os�8҃c�U�G���6��a��\�H��1�"�y�d�f�0_(��IcA�,]ojն�g+Mk�>��p;��9�]��W_Uq��n��I�G�7y>A����������	���Fp@z&HtL�H2�|���C�
����N"҇�-��'$�<�V�9:�?��X�*ząo�;&�s�	\��Y�!�`'@oȍ����! /��`�w�R)h����2J���e/���N�N-�g�$|�7�b��eK5�]�!�W��Wj0'D7T�r2����H
~#�B/��G�J�=ճ�-˛��W����lJ�����}B�	*�G���fHp'�T�Gg�1>q2
���~��p
"w�A�8�j�b�wjI���N���g�:��q�e�]f��ղ����%�
����g\�l��N��3���6!^�Zμ�>j�B�D���������{��1*�`��WQ�+u�wcd}rI�5��Ka�:��UD/1�0�+]f��*��)�GY���74ɍ ���Q�0R�S1��jKH2I�����{�y�	8xC����_q���$���]���M�d2 �e�&�0���8����a����
��i���b��0IY���ϡv����P��Y����'���h�%I������i��X���x)���?�=�7A}R<D��ؓ]��(�I،AW#� S�����tj�aBv�l�,'n(_�M�:/�1�'6F}<�}����p \�i���tA�F(����,O����
����/�
Qo;�1
>��	�[yɉ��+P�9�$�����~�Ho7wg�u����g�S��K�o���JK�r��$w]9����G&uB�Ǚ��8�s2�vW��'-l@~���&�ꪛVP���i�'`�u�#��y�yr,JW*qm."�Su����"7���ë�#Y�u_����Da%�z��ڪ�T��/�\fd)���:���M=f�Xv4�tp�DE����ʹ���J���2�%���q�
ï%��F#��lm?b�C���KD�|�R�"���Jڠ�~dD������~��X{ Q*$�IA�����Z�0������a#��7��\����u<�z�u� ��CȁN>=
i:��\�4c#'�8�6�pV��,[痜/�Pf�-��P��Ӌ|�q��a�m��Y��![�R�D-
�
E��b��"��W�m�8[����l"2Q��nr�F�?�+M�e'���ku�eHf����9�\��}I��E�"X��M�F� +�Y�23���4Х��\#��Lݖ��$��#�KU&�E~p�EÇ	��2-Dq���瘑;[�Ķ�s��1O�t]`=e�b��F�x����挞@��nih��\8�����'�"1�H8��*�W��\y�78jD/޷׽(�R%�y,��޳!~�X�� ��~�����p'��3�Ţ���F�*�pe�W��N����z���-ݙw$�zz:Or�F���	*������H.h�ʍ��!��z��Go40:�`�<X͜	���*��KJ���w;�Xt����"@X��~�����J�{7�l��g�@�p�����!˯Q�	���m2��"6.�����|��lx��Ƀ, &���b��\�E\�l����'��Y���[��oق-��Qa�߱��SE'TT����DD�	��p��H+����o�۞�t�4YO�ɠ~��7N�c�GOt2a�f&F㳬)SC�$�2?���=&���^��`�LS�Tu��y�|�z������1���`dڨ-��{�=;1���-��XR�~�LD�ԩ����������X��"��=�p�O���c�3b�g�k2�=�:��2��ZjXS����CL���d�[�:���g*q�V;�?[���.�¦��H7k�d+�,X�c0P!�0	`�1�z�ӵ��c�6`��9�dǪ��x]���$�s��j�9�-�di�J"��(�+E1��_��m�F`�$�1��:��3�Av� ��}A��hxmA|���#��I+}�1�� j_�߮8JZ�Ϡ��S�Ê���nH6���W.٠ځ�Û�)�QS��Ƒ2�a�F�,@Nn��(l�^%J["�X�P�9&�n�q/D�*�VJ�='0��������Ai�̿�m)���O��^��@�db�CS�X����=lM�n��o��Yէ��BxNv�$˒+$Z� <�5���S�"6i�;��⣢vdҔ��(w@�'u�>�6��_�Q0Ϧȵ��4LV(]�(�hH?��/Q+�@e���}�d	1&s�.�ˀa//ҷd&j�I!^���҇��c9Ju�2�/��)s��%�����M�$ ���k�5���!ڒ���տ����`oG羈���3%��+@6��z�Z�h8��ߍ�&�����T�ˈ���r�M,-��B
��U�O��ެP*�_h��n����R�|�r��*�4^�텲����ꨔ�@��O߾|2ͅA���#�W�}^Μ�w{м���� 1{�!��{�W�����AL2my������)�5�8����!�[f<�����ʠM����e��2�Ds�w��&�Ʌ�Д�}��9;��uH)��o0���ޯ�.I�uz;-�Z�y:�DG�x���iw�s�@�[cg�H�El!/ �b����d�1��B�3����/>t�^�����Ѷ�3M"�|6��MNwВ�m���M`b�CҎ��h%F	_��dj ɥ����8U��z����eU��|b|t{�^^ʷ�˺x�+cc��:'1�x[e"7c�����2�{i��h����k��I�1�z�B�<�t�J]�OO�ְ�H��w�>Pu�l7^��� ;�6�42X}v�@e��w<ĝ�㓩�p� pq��Dڃ����m��ƶ%�0�ء�i2�t��ՕEq�O��LC�"&�$/� e����j�^D�iONZ���M5jBb#{�`$����k,����Dsئ��\ː�t3�L�¼�t��IAA�p|��r���\d�y��K��>'8�fYe�^>A�nܫr L��T�7�>J�s�R�7��<t����|��De�s�2����t�VW���QV��Z*����ڨ]0�O�EP�,F�ɰ��z�����JS监�˂������O=��qi*���f�O�,#�R��%g���úQ϶��-�����zA���� �(*��v�Y�!����C����;u��G��|xL�K�-�\��_�k�}���+���r(9\4�٠�ӈ���a��w+�{���2�g �G�lP�vO�6����IH��H]sY�����1kb��}_��8mfMP0���w�El�vl� z%������	�̠H\��3�.)~�s��$_�ҿ�	�:qf;6͋;�	ŋ�`h(�%�u��Y���%p��k����0�=�m�O[�A~�I7C�H��"ͣda{�h��^������F^^J�Ff�cZ��]!0�B�lG8�kye�(`{쇹@�FqP �����^� �,�<1q��ХҰDē��2���OX��1����n鐘0�I�q���v��n�U��� ���
�4C �^P�Ϋf��0Z�B�UY|��MK5{��A����r-ϨSB��;�
TBkM?�B�K塸�]��b����M�)@Yn��7��X�#����ф(��G?;�y�OKDw��^��2#��p�hY�M�A����h�(�b~J�QĖ��mb���<�Z$QP:�йv�~|��`�
Z0l��-���p��֦�:�*ؽGk��p��-� LLjCz����Z�?�DB��y9Ǣ�2�{�� �l��h�"�{��E}�3GIԻ'ظj&������ W���wi�^�7�g-USS����J��琧��='�Z��
�Ó�P~�o�Y�>�n��n�Ơ�
��gR��hg���2�x���B�FCZ��C=4��7�$�\P��V'���ap�@~ҩ���8�7;����#�̣"=��+͍�Ku틻?��'o�t�:��u���mȐ0�I�̵J�U�7���������^2I�x�����n|}lY~���*g�x�56��έ����5��q���)v���[�o���ܔ�Gǰ \_�!��F_k�@	�*2�ir���c*wd��:��㾁��	�xt��0B��g%�VVݨW��*�2UhXh�s>.$w���.
Ɗ����:Rshf�|\N������)�ŧ0�A����W�DU٫E��lp�j�����
��'��p����B���]Ḓ�Ԫjѽ��د��q�� d� @q��xTѦ��`S���n��ʾ �*���$�^���Q32�����kY�
����������'���/=p���`Zr2�=	Ѻ��m����P L�N�ǝ����#��Gh7�|���|�;��+> �i2�It"gXxϘ���Z �� 6M�Y%l����!'�"���S��Y��q$9���Q�������B9P�i���I"�j~��-*���������%0oKsL*�y$�fYJ��Ɔ��#mN�x���g"Œ��L�(��ǣ����P�R�rR��J�V�t�u �-��v��>��$�L ���a���ضwGK��rel�a�=�������h��g,U�� @Ϲ��a�%;�9�X.�E�h%���%n�����4=�b��w�ܷx���وIhGTU:y�>����Z���qu>�*B��@�J������'n��G�g�Lcn�2�8�kV�Fզ'�O9�M0>�� ��K��zl��h��"Y���+��Q�z�Z�^-u������w����}+\cXj������7q��Ɇ4}��CP���>���5�7�#%\6w߻�-$�mr|�<:����S��-��`���ߙJ(|+4�r����>����ļf�;n����'�R�����,��a����E>�Rfz�v��)7����ȉw΄���(����Pn����H�o#�1`�ޥ��g���\�۵]�Z���L��*{�#<23��>���Bc�k/a2x57���8�TO�7�e��v��X�qt������N�$wC�!��!f�8��C̒�o�Eq��0ZU$	z<�o�åi�M���I�Y=?,�s�^����ZΨ�_v⻣��z��i�ɀ�)���&#�,������ڎ��{�W�t!�I9e�s��5õ��
�Z�F��v��@��_+.F�� 2���!#�SNj�n�U�D�clZ�1qG�]/���0�g�t�;�7����@���:dq�ғ�k�*vKO�E�yAP���BY�?�7��ش*yx>X��Z��^�pbk�Eۙ<%!�@*����]����p	�[����%*'�B�&���h�ڱi���?���{-��!Q��*د�0X�\7�҉�YV�3���0�>r.����D7��u��Wy���Q4�s�����+/�u��:Q<�rx���Oǚ�Q�X'��;�L�̦$
2��\Qy:a���NusG���?��.}��қ�s�Z<_s�����)	ΫF:�O�pC�::����n�W��ðJ2�`��4��H�k.GҜ4z<�n�8s��R8�#�퉢��ȇ\9Xn�0|1���N�!�곆�ע�#��Tw�--K�r�Y�u-Rt�j������@,�����pk���<DZꬒ�R���t�pż	6X��4k�.�l�_�tU���[+%�#LOiw�2�V?P:d$ď/�{l����
{�~J["3%�y����O9��e+]�[���x���=���]?�[9�'=�,qͣ�����4��z��~�N-�k��z�;�d��0�!b�ῷ�[Hr���[��P?��+�x��������<l2�l�F �PQO�� t_-����E8��}Ɇ�@�M�d��-��J�c�]Iu�%詉;nѻ�)����Vg}��jGB��'�N�#�m�0��ɖTś�
����O��#�:�W\��YG��~��[�f�<��J��^�wL�4x��=��!���T��Y��9�������12B,���?�e�!����jQ��	͘��,�iqsqV?�>t�A�u�L�������F���F�V�����Nz��G����\̢}�h�s�l��$�N���3+/#��9���D')Q//p��E�V��E�Uj��hք"@�V�N�a]Q�)E�ɸ�O��� �f�}L����.�:��̌���n+=3�6��u���fW�~iux0۹D�s�/�~e\#�*�e1��'{� ���$Yi@t��)<��I���9mv`��7
1��<:,�vhl��e ޴�����~xA�KAPoh+��Y���\���ń���w<�!��8e�K�3�ȁ��]�{}tܹՁ���d����mp��y�r jf򴂺��i��u�4���=�Y5滎�d�De�\Zu�y��S,�*����@�~5�h�R���z�;������'�k��ɟVY֧�a7����ۈ�� ��G(��C�|v4Y� ��j�q땵�iK �ʓ�l]�fq���1�P@*�xs] �L�f>��11��<�B�COY��?j��)�Pa����`�F�	�C49=�V�[�;��^�vx�:_�>����]�^��^�(���h�T��pˊ'���]�{/:���^�$��sM0�N��8�{�X[͒*��?�i**��"=�b���(W��-�c����\��1#�ٯ �v0 �6��!��a�>z�4˽���A�9�Ǌ/�{�X��Y�F-V�u�z�p��M���p����;D3(�pûs�����Q,8�b/���fD��I���z
����TЮ�$.Z>��}�0�F�b���#97�}?1���r�MĄ��7��W�%��"#�e4���ꊑ��Dy��m
=/lN�u��an)���"O�+���7��(^�Z^���ڡа��zF,f�7k��SgP\*��0�{
u������]2��u�B�w1�}Nή�ڧ�VD��n"W���W�����zsf�*ߗ4z��';�6IE�m=	����A�k�.	�r-[�?�[�" �֒��Xl���ǽ����p9�p��z1bd$9�L�ɩ<�td�۱�mY����������:��XP:����r�<�d��^�	u{���"mh�R�{νq�e�Lϩ�k�O�ޏ�3.��mpr��ݟ���NB��o�4��� �6y��/m �ka�F��ѭ?j�ɶ �`��+�C>4}'�:5��.:����ς�[d��p�6��#4%�9 ���+4�g֯�.ftܨĢ����� ���\v�����vY.�F�����"�vu�[�S��"��@:�ɿǫ;��M�=]�c�z�BJf־�� "��=��82;�/|��]�{w�ji#�^��SY
D�D�X�;����PfXn!����c���f��H�ne�-�t"�ٞ��k%´�� j�i�f�I �G��3�T������v�|=�¬�C��F�!�a���Ozox�P�=J$\5C��z�W���Y��
��8��}8tXc弞܋�]ݞ�[Π��T$]G��(-�e/V�Fd�2৽��%+��½<ȓN�Y��6�R�b�7�7��U�BPe�����)���N�9�=��'�͵��ͤba�7;i�zn;��k/C�QbS%Ը��[p�D�e.4���vij�V��|l B�İ�P�U�&�m�����[�y����~�#�MX,K��~L{���E�Q����^^K�� �4��hǮ��-��Y��J�ed6���8�
����e,��m,���-r��Afn6n����*���w��,G��d�/��)J僽��Ihpܲ��$�h��� -�>-\�����QG����l���z��"W��lޅԖq�bU���k�'��h�m�fnU�[J����6V�b��p��T.����nZ�KM�t�@�o�jY�ˎ�Q�o!Ȁ^������17���#n���Cw�i�Ž`0�6<��%�W����N��� I��|�Ш|pH�J� �`�с�Z�/F_9v�co�G���1��;Z�7|㭥G���i���܊�>p@-ϟa��9 �io�E�����v��oO�e�!z�[��ՉצQL����"��l��.�∅2B�xU����)�[y�ct�;@�Jv������+���1�3�2��]A�"2�YT�ą}��)F|�x!�1�k�+�pW���p��S������"2���F�hK;��[����ƣZj�M1�$y��'�sli:໪�TF���2`��=j��I<1�"���4'1��m2�x�GJ�+����3����GJe��B՝�C�iɎ��Yކ�	����c'�vcll�^�ar�|4E��?ڤB�뛗��sf�u a�o�������v\�%SXP��y��VbŤ8�ha
('�Ub���52�W���
�{׫¹���ST����el�+������� H%��<�8/��k6a��:4 O�ݜ��HZ�L�w���.�}jA(ǹ{�8�2M�Τ����v�kb��R��ʹ��H�6p����
z_[������f*�ڗak;��ۅnK4u%(;������"�!ќ2=�[}�Kҝ�r��C�q0qԻ���J��A���2��A�)6I+��l����{�M@�h1zː��ޜ��c�oCĘ�?hgy=����H1%�.��g�P�M��Z ��a?�[b�JrȹH\� iz	�VYJ����xJE�1��`'N��3u$����Uf�ڰ�H���<K�rtڸV�֟���bұ]HHLТ[,0�&��M��o�'+#�b����j�qBu�K����d
��