��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^T��Y�(�,Rx�s{\���	����jՏ�z��7�1��k��y"-��r�VO��������Ԯ[�;�2w���*����r���$�}�����OC�޲��D���,����ug��)� 2l���˲_�`!񘙿͝�N��N�-��^�k���o
҂kbՄJd���Z3��<�`
�������%��ٚ�=��=gױ�Co>���͇��k��M�i���P!�G���jEFВuy�*�6r
�>ǉ����A��M�w�zHM��������[�y�u���U����q��;,\&1��wX�4jv5����hl��~tSCP3Mw֊*�C��#[��c��6��3�Xw��b^�����c{��TW��X3Ӣ��D����!����� -;���6�-ȵl��a�uCP�PL֩8�@���*��^��PI��s*����hG鼆����W�O\��>�#E8$4>W*��5����EM.�jA%�9��L� ���_3ݒ�x���\�ę�0l�~N�j5C��V��jtfB��Y�3���|b.�:� r�W�컯ܝ/�4v�����ˍZ68�C����y-��~/�e5����/� W�9�7�1��M#3�hM��z+���먾=�k�
�����9���]���������>a���'y��yx��=�>Xa�'bRcx{�9$��P���c��n@�oq{���|�����@iJ���������5��}��X|������[��=d5��#6����U���0�Y��&G�:�Z���Ai����,1��M`�8T�!z�l[�b�T�>��qF���01���X0�MX�ڹz4�_b����_�5��8���W��-��?���������*AkeF�tD��.����k�G��o���%[��`��+R�9|�d�O�|Z�k�j�2Kv�x<�,X��ϋ���j��5nJ]e�o�~z
~�  M-�I�/t{B(*H����M�5'���ڌ�'��t�.��/5Ց��}���1mp%��Q|u�>�����`R&��-��j\����(3)o;�WՑ�f�޶QQU�2���O�Z�%�����J��0~J	��*^���F�b�	F�W��=�} dO�=+"/�y��|#v�"���Ҧz���nT/&ࠪ֘>*P��\�5������VZ[n��'��/`py5#n"�H_�5��N���E���e����U��
�{`��:i�Kj&�Ȫ�
�ǎ�8@|�ʌ������ ��2�7����>�VHD�����.gs� ����X��?�>o���WĠ: ~�AnS�Z~��o��GI�Wã+^9е��=���V[�{w��$��w���,GI�=�m>slrN3G��|�����8��|�.[m6��ӏ�O�׭��������R�w&E�sa�c,F�[|!�3��6U0i��&ŀ��(a���C�Xs���v�������K�����=��0[�@ٜ�:s�6ڕ����W��N�hYN+eXۜ��`�R.8bL��OrGunK�9��h�F�!������dC�Vp��f�O��U���6 L��S����%PҊ�M0a�����e�-��X��0�kϳ�"Hp���:_0X�;�ϓ2���eI�<jɘ���1'�h�������DC'��qy��:��C��6��N�@�����
UB�Y�NY��p�\�1�;D:��p��b<�����6��	�nZ1��tKD��W������)�*�qp��ǢdQH��K�m�Lx������Ry�v�"���sjɥ�������ћh�0-��ۺߕ�A�#�H�����c�eH��'~��N0�bȢ�.�gx�"�u�����#O�g�����ߴױ����8����Q�.,Ŏ��(�&����Y�s�au�s�S����	%���}���LO<�����V�$�z�z�[F��e�r�O"������S�_�^6��C�o(�;���VSB�/���%V�>��',�P3*��y�,e�)�ψ�q};��s��$P;�0Y�Q?#fLV�X�����潄��D^�Qi#���:Ӛ��`؎?:H�#�k�;$��	��]��sIO$	݉���%�U�f9<��y��(���%�_�%�3����Q�u|�*9���h�f��j�����e�O��"���n8\A$��~�F��v���2��X@�[�`[0Ej
:�� 8��șN�826�0���E�Ga�Z@��̳��C2zYǠ�wUcS�QW�˦b���"�P�$�}:̼�W�g�7��9�����X���n�ſ������G�����j�^3[��zμDP��	��Y�a�ђ���>�ƍ�{���/Ŧ7_�V���;uyh#�sc�2iҫ�~�&�l=	��\D���d��⿞����Ӱ����w��f`�)(�wԼ�փ��8��� ZjD�#�����HfӸ��$��d0v�@�VsV\��
O�lnU�c�]����Cu!_����RF�g,`S,s��Rp�~Wd@�6��n��?@:�̖e�<�Ji�$#��
�%oKn��RB�A�_T�o|�յD�E�0l^��R$чԼ96�����������Űxכ��* �ND��B�N$K;��5\da�,� BO���#��*f�|�q}H�5��ٔ��J����4�Ay$Փv������?�ÍaY �������q��!+�$������&��"�#Te%*u�)cG�Y�h·/�c��>[��s��Vv�8���,�,]�=q^;"wʙ�zϢ��{웂�e��9*���r,�t�su��͓����TU8���x�$���\�I��	�'�>���\�n�6LL�|t���Dbʹ�����O?-�{���P�gw�|k�����2r\m�ί�t�������B��Ӗp�d���W��MV�m@F�?��r����d����zb��]b{���cB�=:[ծ��M5hކʑ۽a���~G�e�ay�XɈ�I!��Szk���F��R���0�G(H�{�X�Dm'�����}CAZ�Y~f u�!D�Y�z
��))��OXk��A���3 a.�@�INnX���f���d�a����Ҿׇ��~q�S�ǥ���qX��������w����6����w��5,(e���7׆�,�ũ�"��I��+�F�M�0A���!�&�.��ɾ��c8p�/�����+��>�u�q�%��̭�G�������NŒ��b�k}}���g�0��͔X��v6�Z���4����숫����#w��"�%GD��zTj��[ʑ:�Y�#�Y�*�]V+Fr�	��:�;�6<�W�6<#��%�	��~�z�G'&��I�}�_�����>h��!EQ6�L�;����̂v�m�k�j�1�r��ϴ%sCa��߲�^���F����[���4n
Rs ~���j^	�ON84^dSQ/��j��]h�P~B���L2�N���P]�v�pE�Rb20�K�H�"m��`=h[��-������~lh(�����w�m�ڇ\i�81��P����ϭBD�P������}E
� ���
�`���v�1�y�sB �$��!��X����܂��
e+'�}����,[�ѝ�

���*���	}�r�[ 	��m��h3��R�v7-�_Eo��m�+�UO(�P���N�X���( �o4�]�����W��w��E��u�3L�n���6��;��|ū��U�u29�m)9`K�O�K*�_���e�z���Y&��Ёu�)``�x6F��ҕ�{�`�v|��j\3�涋�@������*�Hmϭ�u����s���_Y��7��g�����|k�0�S��k/�)���z���S�3l��h�	����A�1��j��b��
�?�D�>�����I�<&��&��o��/���ю���N~�RD:���+�P��#V��aAS�S"ل���f!�fƲ������:D����I����6װ�C#0ku}�E4�"<e7�$�&�3�텛��V�����+9+Pq�&v�8��"�:�J�$�br�O��n1�C
@,�Ϗ�4Yְ��`v1i�.�3�!�qA�G
��j�3TG����1����_�u���CvuQ�xi&�0�o�_&^a_��e���2*����5�p�l����)NS �@dY�\S�ʀ���y�Z��j�
w&��A�ntO߰���>�d�����ߨO��E&+%o��0z����u�+�n@�j�av�qwLM�9��������(\^o	�4*U�H�A�.��2-a_9�k���?*j��[ef}�T���G���n5d]�سE�{Q����f�_R��}�hR��x�E,�l63ĝ�,u��+�`��q�u�y�4���E]c��My��1��(jۀ˚GvE�&D��]U��`[�u�W�3`D�iaqV4���	�~x�eDq푧U��<�3������O/�~����CUފ���%��#�����Ե�,��:�8k�u0I�&K�]~����1�X�k3�s��~�4+�m��;n�	�S�UK�Ĥ��S�
AK{.�U�2�(��w�Ҍ;eH��1I�:ns!�x���*��l�h��
��hs�l)�:�tfXM��V%��r�xfVO�K��
R!�ab�2G���^B'^WVS��̗{�̄DN�:��Ɂ��~Fb@�`����<
!�R"SH1(ژ�4Xyxh��e��.�y�|�;�o0���d��9�`uW�rp�Z���2��u@�W�֬XX�zim��i~Q��-M��֞j�'����4��90y���[��s�mb�Io�+[UB?(bs8B	b3���7)�N� 	�Q�Qh��߆���c��li�;�A��2d?Q �50_5��P�tͮ|���%N��>_��)vy��c�&Iw!nI�8��
�m8���H�)��:���-ޙԵ�4������(:͡msIe�̔`������@��]���B��{^/��Ce���������ބ̱���w(Sd�6�'.W_��� -\�V�p�7aH�:�#��]���R�B��YZ��b�v�Ժ�<����-����k��SM1~*��S�Xw��lq��F:���=D��z
����!B��m��t�Qc�&9�֕�(,�0��qX�H���1��;�?p$�O�O��k|�R�� �V�9!��a��[$��Wy�9ew�sP5Lu���i^ԂX_*�3�ik�zQ`��;��"���q&�!��d/奼D��{��3���g_����t	�B�����p�~�وc�`�EW�����aQ~1��ޞ!���κ��p��$�HSH�u�������mv(\����5���f�~�u`�����;�W=_��,������*�V�վ=�@�#W���ɱ�9Ə|�b5�:�0iW���Z�X�j��Q��(s�O�w>�gJ��4T7a9>��SӄA� ����6R�h����Π�tw��D�����i�}�Dplu�>_@��[CZۇ���2��\;�5@���d��Z��ruu�ʁ�,2��B��v���I�:��+���j|���I��=GLH3A&�a0U���-�Պp��RB9^�h����n�,�c��A�������)�~�u��֊ Z��L]--��b!�ʖ�^Xئ�2�>Uꦱ�V9�4m%�n|�,�(Ar��@��Q[�H	���Fc�!��jwz
�=��3�ט�?�w�d�N���Ȁ���DR��JV`��;,lA��\�^�o\�R��&�[��W+��,ݸP�g���X����W��gr��S�$��h�.ng�c�L�zy=���*b���r��?hD^�ǯwǮi=ꢷyp��7��ot��},�!�Z�Ȕ�wS��*a����EG��4�cC+�a3�M"���pxe!�0�]�8R��r*�.x0�M�*7p�4���3�˥��@]��Ѝ�Q!���Y����o�`|�慜2~'H��#�}(���0�a�Z��`ԩ��d��x,����	���⬏�5�:7��ie?IQ�}K[T ������%i��Zʨ�n>�^�p�I��Z�]�va�,��zx��*� QJ�vԌa_F�Cs'���m��BAN�T2������S��%��{�A�b�/@���K	k�gӳE�Ŕ�l�-�0��=e���H@�Q��
�W��a�����E��l��Ou]/E\�̝�PZE�7���5�hI�~��I���p7�Cj�C�����FFǜ�,w^i�V�(��y<,;s����Y֒M����!��O_�t�6���GH|uc3����[E:��ҷ�ш�IxYa�)" cxg��"z��\�.�g��fT���;��>V�Da[yZ /�d����y�9{j��e ^�-��Z����*����k\��9$d�[�@FY��抱�V�Y���Ğ�e'Ҋ��H2�:M�
7�kB�7����/�>�k�ac6�D0J�u����5&s�ᶟP���F1�?�z�,X���e������[��j�Q�b,��|��D��Y�~�rWWN�:2��҈qXv�7+oE�`t^s�8��2�<���	6b�m�8Ƅ�"�m&�Ə�՛?i�.��U������Y�����]��mG��a�i���2�������9]��icdն@vLp��F�G�50b*���!aʪ�N�֤ �+i���EK�h�����}����:���yم�c.h�p_!_ki�t��9���{�~΄h���H�a��ݕr���[�>_Ü���v{W*j�f�4aNbf�T)o��!n�H�e�f��g��{[|O��5���
�(����O�4 �N+�R�'�ķ�d
�!O���- U��rƧ^+�R��,���P�d�0��i �{�:;��IG	D���q��ᮉ�����������C�G�5bR�EZ^�Zx���:��?��n�=��lV�Zrp�s>/F��R&����.p_�>�A����?��˄�i�e.M˯rH�g��>�����* ۫�,���U�.����?�;bf���
R�^,��U��N/��y�jP�v���X�\N��#m���;d�CDP���ȡ��..**_�_���'��껖���9�vL��`A`~4.�E�|;��a�a��[�����:��1g�+B5���{���u�×�S+9�H��}�n���k��X�b%�Oܲ�f^��@��@����R|�Q?@^��� �-�_��y���t���nw=o觚L�1���x 4�H�QC�ӽ�J⏧o~D7�f���]��V�T��d���=
���I��On.\?ߙr��A������{���c,+��\*.��\�p���=�DԬw�ӧՁ��<ҫ{�0l#G Ԡ"���OIC~��B�i����k!鶕�dOAc܇c 7�U��/& ���&_���7�#fMRE�"0D������VY�Q���.���	�o��,�J'�U�w�v���++oDC�f����B�j%�2�
������ؽ�խ�WGUj��q��a����l���N�*H|4G �+W�%�~UW3�F��j�S.,n�Ĉ�0= ̫��O�w
V]�R�o�5���h�c<y�Om<��ж���F��[DG�7�M2��%�
<Q��� ����N��Xͷ�
��u���b�&��}�ǿ~�X�h��"
�4�������$��{8�K�U��u_^�r��f�$J=��H�Z�	��M�f���P���1���dg!N���}�z�j�Z���R��k���ģCd���X${��)N2@��85��آ�x U������W`��C<)��"�ޚ�ȩ���h�"�eS�\-(:hSR�&�(�^L����
��h��ZO�w���!���3ğu�3�#�uz~�.���#�+�FD:2��,Y�bj�a�=S�X~�h�F�^�u9r��ı�|�!60�͠����{$^1��6�xS�	H2�B09 /~��+�g�kr����!��X��8-�r�U���*�n��M��]���(���k�����;{0�m�E�I��W����,����?�7}P�m�4�]���}}�<<�|9�Ov�S���Ӝ��$-��ƕ�����uE��;�?X�r��4�J\��͡��cJZR��4CO�e�j:�lHw- x�N%zs�}U����o]��|��7[���kAM�ۭmL���u��O�@�2��7q��Li�o�[qA��w8��a��Qq���� .�]���*D0U����(�B�(թ�,s	3�={}���������g�x	�%̴klGx�a�{�+wm	��x��0�_��;�OA�\Y�,�a@�j;a��c���#y��������
��+H��ׄ(Ixb��f��u!������4� ~��?��	ND#!,�L�	���.�����=@_�(cI�;)�L���|����zV@ˎ���B��o=
'u�jT��X��enc����Ђڼ�b����&|h��Y���-��1�vW�7#'Zv��>TϏ��a�H��J��w[��3EL����jҼ_<����\U��]�/���J�I��oE*���`�&d�p	��L��RO7�����~����|���	/��H�\�>x�t�bZ&Z �����}��T��<eK�K���9M����3�F9�W��}`J�tKt���J���˯��K(����u�oa��L@Xg/�I�j��2D�^��⺗�bй��}���.�:d� Z��9~�WK8��A�Qk���Y�uͭ�ˑ7Ջ���E�1�݅g>+X6��u��\��a"e��Ҫ>��a����}Q��䲎�[Lw?��|.7^(��\���Z!ynK����<��[''�~�+d��~��C�C+4օ�RCb�91���B�tz}��+�J\�n�lq���Ŀ�lS1#�VR�W��u{फ़�z�)�}�q��__>��aqiHH|(�T �O �YպZ�)b!b�-l;Ș��LM� �6��L}&c77*�ÝŃ����QE�NĿ��?>�.�n����t�� ���ME�J:Ҍ6/��H����MݗV3�+ʻ���#�ٶ��̩�{(����>��*Y'6�i]/ (0zc�8�X�˜x�O�'�.?K'p��K���X�#^C!kr�ޗQ�m_6���;��HN�����{"��ވ�Ww���n�D/$���/���8vx��&��7#�M���&ƾb�"���ZMg��f�u �#\�^f���=7�ޏ�do�6t;�����%�+S�f6/���Y��dDB�k����^����J�Bճ����c�+S,A�{J��הpEŗ�~�=p��u�p�jȎ���1�ͱ&Y?k�n�8�vq�E��
�;��5�̤]��_�ؕ�:�kT識r��{�i;���P(E�֊|..�}�hd���n���_��Պ7N������f�GCo���|��R�-��d&�_��Ye'(�<:�z\rh�� ����B�I�D~�C@qє�tF\<�5�E�-�V�)�\�&��O6�H��ӊ��i�3U 6��_��a���с��t�]s���w�CtX
��jRkӭ�L*}n�ʄ��Z\��kTɚCg�?��LRX5m���2\�S#.���%w��:+����wKB_gL�~�u�����d���t'�jӪ��nZ�@�����}��{�k�o�.,%��	\
J�i��*�@yr��p4�6o�/��k�H��������e%ݺ�� ��?6P���>,��C�o�=���@=�5f|x&ByT�;�&w ��o�̴��"���Z��3�Y�?
�a~M���,�-C��-�̷�����<��`�f�h�'j�-}#'�B�9�ZoGѽ����|���Ete���pӛ
�c<�mEvmN�G ,§2�1Pdu� ��A]U<�r<+o�K�
0 ����2\��Ͼ�:H��ǆ���{������q#`R�<��+V�o�]a���l����	����v� ���ɩxr����&���GX����d=�,I�ǻ ��`��Ң�.�����K?�X]���$���Ю��̉[�qgH1PE�����d���Tg��ޏ���=z����jg�S�V���tc���� ;2*1
?&h��=�cN��k��
�����e=����PQ�Ǡ��3a���Ϻ��+8���	��][�iƄ�ϣ�����̔J���hA����*��/h���,�.xR���������Y����qC7@7 ������@j��Ȑ/J��<ۿ[qΓ�}�35�sQ�݃�����,�(K�U)۾��_������c��ܡ;��Z�N��2Q-{5��f���%�ٸ���l��m��v���7���J����x�`�M2l�?6�,D![��g�HmN��TE#-��^NK���z�TS�I���9n����H�_� ]վ̏�
��5�ó\���Q�b�%i��|�S��r׳�x��K��Ǥ��8|���~Y+��y>{�9 ь�",]�lh^y'��!�t�t�d����I���NR�L�;�=�qڍ��z��nH�֌ �ȫ?V��,t�ȡ<��z ����|��c�䐄:4Fݗ��0	
���摺�Ǧv���UgO���.����[V@ߨ^�� �a�h1�r�6_)�;�0���.K_X�.�_����V)�T~+����JF3��r�=�"p�$��=���U0����:P���<���.m�E�)�[�����Izh_��㞔 ����vͦ���&#�Ճ�����wgP�-���k��`��h�l�N������ ~��ً��̝J��p��{JB�怗qck����% !��0�O���[�������F����u�B��Q�~ax���0�Ykhʋ��QX��}\����*2�FcQ�	!��=ٴ6ժ�^�կ�p���XI%?��<���7����o.iz����EH��X��Ät#v���X�x�o���s�jW���,���1T&د*�p��j���ڹ�b�|�V��7 B� -8-[#_]A�Kݴ������M��R�}N뷣�4H\�J�̩ӂ���o����%�ҋ��p�4������tt��{���;hN(�j�dXl�f[��_�f����2;&��֨_���o[����%@�Nf�n��Բ訚g��B-�+����Y3�X�����X�ny����c5օ �m�bh��T�񀩂��!|�������[zg̎�8�n�
�c�3?��2�+���w#0Z���>
����Z���h�<�i^`��b��BP�څ�1��l�nY��a�<�ԋ���s��T�j��7څ�]�)���b�~l��IF?|rI�r�R7�����߰Xg>��b���"�X�������<�Y�Xj����?��>�A�*����NpW�{�=��G���F6��cSxU��Q��r�k"cOvP5����N��P�	n��J��{
�L��	ߒ����F��TY��\����1(�>����bv2��������[U8�a	��lfK5�7&�T��&�l;o%�g���O��>�{S6���`�E�t�Ӂ�TvEJ�]x[�b`��Y7�qr����EW�%�8�H�@�ųԸ���M����3�������
����ͺ�J�oj)�شt#g� �$�H�6v�����\���^�����m�	k�9�!/X�6+�"R#�+\�����r��i��K���xt�n�SG�!�:�@���+I�(��c_ܤJ���3��:�u�Z��Ĩ�ݦ3�[@��&!�Xj��2�KΉJ�S+;��m$�q0�����pW�ǖħ_uod��v�>�Z�$��V[���Z|�6<da�S��)��r����J�����x\���SZn~��,m#�7�S�<�Sqz��׎�i����䳄��Q+��Nv�"��|l�����ׯD赜�����[ƪ�˒jy�����duh{��"Fe���Us����Csd��򛽿@z����A��Q�J�^/�}/������v�|쥖��q��2����^����(�����k;Hx@U��������c����<�Y[��}K���;:�U<�݂PZ���;t�ЖTk�oֽ�A��
�n�=��NN�N���9�D��/M~<�l88$(�dt�[5�&[R�~Dg �xޠ,-������a������o6�9d�L+�ss���ŗwkh��_et���N�{�;]n�����蘄h`R��@3b�<ɉ{���F�i�I�ߓ���w��I�.∝C��lޕxX�S)�C�����U|T�v5��P �$Ԍ�bA�=k%E�`�T��C֚8dU�-L��kr��-X1��PV,����z��P{��e���	��5
�}�wœ�����@e(+܇��U"-��ɘ5�7�v��(;w��B�����E��g�-d!�6��e�^��o�D�iq����/:V���x0�qߍ���.���?��'rx��-巜0��@zkjUY�h����������퉮y=^��>���ڎ��y��VڅY44��p�[9(����%c8��N�FּV���V�:ط�<�Z�U����7;�4 NJ�f5�CSe�B�oc��V��ګ��������.MuX���?2\�q`���B:+�ϸ5����{���[j4C���r�Ȏ@w���(�e*�/���UኛJ]�����^���J\��	�#���(���
����S��0�1�jKn={�`��P���\��	����8:~q��(��b�i�uC_�y��;���q���=G�Q�3ؙ�cEtFQ����7&���neZ��������n�	:H<mM9f�@O���J�����	�~���@�{�EJ��	
�\n����Q�z�;��[��9�q�y�	 �0l�y4����L2��]�^{���Ĕ�����;El~��0���L��v*_�k5d����-.�yX\,�
�P�[��&����NvdBߟ	��V��8%�R�lĂ�q��]��̥�l���1���D>�!�s|a~;1��^�����*�;�5�9�pV��m���c�CS�h,<<���{k�}(+D��$e�d��>� �� ��K��&��S%8�럓��j�D�W_�����&A$���p��X����_�D�9h=����߼�E��ؙ+�M�.��z��6��wEj�$���Ms�����v�z ��!�"E�,g���c���u��z��˰(9��ђok _n+�WC��WY�5!
8ѭ8h�Ks�d� '�1���_AS[�vI�4�J���H�+���慨C����M�az�\��	< �~�m�"�e��i�snzy ڎg���o�Ja7�.{譡�.����#��)Q�t�GDt�RVF��m���~>������P�� �	�.w�-J=u^�.Ai���_�����nq��bc�-���B�2hc��m(�M��$NQwZ�G}u�E�D:S����E�~�WS�?7�N�y���b��Ė�3馜��s
��CVc�>��d�x����v�r�d
o>잎x^e�>�������������3���W�XY�Y#�?�0.��$\-.E�UT�F1�8#[Z�IP�2�s5yySs��۹g����D"��w��@^�Ђ��͋n����:m�/��.n���ӝ%�Ζ��<�w�N}hۑ(2��26��7��6��8���� �=��n�*����_י�`���:��W�tW�)��(F�'3���@�0��IM� ��X%']�a���2� �،�T���I�/���
���=JKkj���`�#&ʤAW�W�KnR1hu�G��S�BQ�� �)t����C�ѩ���o2�ʿ'�3#��#������HE��sEg����un/l���=�W�1�w=r���Ô�è��w��A*\����؍M�n�I��n�t��M%�L�U�.��NoA{�(*	e6G�_�5CI��]f���ts��p����mg�Fƍ�ƧJj�� ��8p����>� �3��p��cG�jJӌw[zM��T������&�`9&b۟{S}���L�?O�H�P����Y���"3�a����J� >\V�z��t����c�����d�
et���h�m2k{��� ��cڃ�@�=�{�:A��z��_x6~$���ιڠ�L[-~]��� y:<ե�*�K�;��V��r�ފR� �`�2�hD)-t�����1��ZJ8ɕ�@��?Ԙ�,��p��n�6�l˽����?�M^��)F
�Q��	�TŹ����|u��n@�� P�;j�o��E�+�/0ɋh�D��q�Y����l�-
���<�l`��2�$���i�+��8!����f9��;��o^8�,`�o���i̥�&ڇ�`m$��l��uq�zZ)	hOwv��MC.P�����)����{��!@�%2դcm�R�Q�u����M� )�,�e�E2T������¬ׄ��H����i+���Θ�>�A��/r�R���'�XӶg�q�(W��?�1��q�i��BF� c?��o6�j�{G��tAg�<#=�]8`�}������chԘ��qBfm��Oܝ��_���*$R��|������ơ�
���+��7U��(��MÍs��ɋ�ڏ���x�Ӟ�#��F�28	z��#�����B�Ȯ>��2Z��Ga�h�X5}���wvL�*�G�nsۃq�L���eC(�}OT#ߴ0ȶ�S{o�MU#�O;�gm�X�����`H��Za�V)���9����%w��$��7��:EUb��wȓ�r��~����O����G����/�����`����>p-���n�l��^A|��m�)rP���y��@���qd��I���c�xt ��n [:�ԣ��]��Ŷʐ���,>�L�b�Q4.i���sG�^y������}'��B_�a�E���W��<�)�$�b���v�$�����+9C@���RMA|~hV=�6��<�n�%���.�6��7�6\>�N>Ґo%_�~O í�9���b�XKRs(޶�M+�<�>��/TW�C6�<��f��<~{��[��6���F$]�B*��N�z~���T�|a��` X�h�U�/��e2��l�Qi��Q��;�~H��YN>������m�����"�(*�\��Ep�@���?�wwK�y�n�}v�ć�|�/<�x	���n.�o��^�8��h��n{'�q���b3���K�ױmO���m�D�.h�F9c�\��V���	�!�}I�{
g
�r���@`�Z7&�Ui�%��뜷�QO��~��I��T_ʝ���v
���/ksUg����zkx�2�yv���&��i�z�('������QD1��n�)�D�]�]���&j
�ށ���]}%y��ږ%�I��0��Ki��_��!��䑖�/)�{��"C�P��p���PnL�}K	��BOU��⺗�ىBZ�g#\,q��b����F�r���%tH靲ף���7����,��9 ��D�[��a �:�HZk1>�H!�=n�V!�_�|��9-b��.Ņ�qY$8��uډ힒 đ~z��BX���>D*LyP���WH�����O�����nPF��-��M��=fJB=)�����́���Pqa�SU5B_����V��n�-�d�����F�t��ъV�w��M����hI�6�`�M\�<�VU����ۍJ�3�-��t
��!��$�r���Q�s��Z'�b����?��8�Q� �#��1����!<�� 쑊W�_f���:z��R;Mr�!*� �^]��3��xZ� ��C����U鶚�q���/~�O�1CZ ;����l��bs�Jq�D�}�s�����[�%'�U)�2�`vt�Ʊ��2�jm����5�����ج����ܾ�����3������OZ�zG�96�6L�%��ii��(k[��GiC�C <�>(b����w+�@�2ܳ��i%49���,��К�&�y%��a��G�1Ė �	FU��Tj�"�ua�'}$'�f�f�$��f��y���;P �Eε;^B�S:��I��N��
f�!�j0�UK��=CU��Q}��y�إ����l�G����u�O��p��RQSa'}��h����ĺe���1w#>��Q�}��5iT�9�����l��yj3�p��6��sW����&~�n&�.�q�.^a4n�W;D���/�k�dt�޽����5&#V�.�:tOӳ��c��r��g%�yYE��#\�i�?0�֚	s
���;U=u������AQè�S#6���E#^��~*�����+�0�-�|m�j����})T�~��I�sA>�p�]��M��o9�H�S;��	�-M���<�X��q_e?cR��dc�!�2#˔�AȪ���s���޻D�}�xu�.����9cl�t�G]/H��������s��hr�N���U�u�tF��x���c0�h^��*���������.ֵ·SQf��`�* at�?���[���0��A
�̀>]�q:k�Fvb�Y�
����Y��zcn�|��b6��N{�g��j�Q�if<���^3o�鬒's)�P�V�����ܝ[�Mhv�݃l�*gĩE.�$'DK��c��la�x@TE� f����/lTJ!s&���A�' f��S��&A���ƿ�J�A{���²t������O�z7e�z������X�'JB�P�***��y	�QBm���F��"�	QD�/�-k�I�l,)��	���B��nW;Ҽ�bP�(KJ��?vej�O�M#ḞII�ec����Z�XU�����q�و�Q���&�|$J;0�ioi�:s��V��J�-�,b|��%����*�T2��]=8h��eI���!�_AM˴> ���`�9$:P�\@D!C�d����ߍ �O���b�]֛�(��Vz����N͕%y:��/`h"_�EO+kQ?}$'+��6R �Ed�89V/ܳ��/#vh��+�WHhN�S���oQ��}�:&紅c�B��:�.HA@�D�t���/K�EvnC�YM�@���}�2�|�W���:R�=>��/���1�ҵle��;�����_x����Fv���lȖ���>�5&�S)I����A�������|܁����&L��U`%3���Y d$��"�^��$�]�>"��_+�W�q��9	:�2�p[�V��-.&��ɯ{���`kN�	�֔Y>�Fu��d���c�и퍔2[j����d�F17y�G�F�y������%��a/6SZocr%��0DSR�"������
$�ڮ6���	S6;Mo�tܠ��Ҟ�[�e�4��D�t`%O��Q�Ҫa���ѱY��яy����� '�����˰�(W��q�,��;�|T ���M<��*��m�p��f�"�MҼ�rèw꘥7Y�E�P��c�B����k���t��9�Њ����v�q7��K,�M�I���3ʝ��H�U�VB���d��zO��ȧ�(U�ؙ���|��(�^< �Y�E��E	���k��F�2�������'��ׯ� �i�i��;�1ҫ&"݄���mӑ;[-�s����1:�f�O,+ �vSSEY��*Zk�1��mto'��+s�v\*�Pi�#��rF�-]֋�Gn�Eu_J����߉��u�"e��M�\C1��eݕ�B>x�
Z|�,��Ť������$c6J����h=�����6l�F����P)�z.���1�y�V�>�Ҁ����o���P!)JĽ��i�%�W�IT=؝�i�t��I\�F3X�����rl5L�^
����%�����$��"�q�F���E�A�fE�QB�<�U9lر�c�lBz�NQ%���Ǟ]��C��?Z��I �o}-�<4���� TR�n�X�g�-5&�͝�aE��L�1�WO:�Ŭ����7I� tţ@}7%��5�]���'�&�,O3�X�KF���3P��[#-���H+�5LH��1�C=�l�*g!��
R������u�.�g-U���&r�k��k6K�7"WB�!�-�1H�^�|W�	2	&|5��^�3^Eo���k�yl,?V�NmH�*� o���z嗑.��n���z!j�J�}���d�] ��n�PD��;���J�t��&��'q�������@�r��FV8�QP�h��.~���*S��5zUmj8�p�!��x]*j�����{R�m���㭅�2Nj5gs�a,6����QC�MJ��/�{L�w���'�W��f�N�~��hxӆ� ��[,�q�AN4yV����u,0�������8�������k�$������2x?���Y��⸿ą5���h���� d\s��X�db��w0���%u�ݷ�*4�]�?��ĺoJb�3߫ʿ7Wj�)b����Iϛ����;���������Ɣ�%�N������п	��3�� ����¦�7[�7�~={��"O��a�38Z[8�l�M�6�n�: �t?��x���g�����<��`�*%��y�te�_yմ9Y5�#����b_��"
�.8����B]����x�m.�m�]�b�yT)y�-;ZLn��/|h�ZSjh���><`m��{�z#���Iл2���ƒ|�q�		���G��WT����H�Wc�[����u��/�6�X�*��n0�Gh)���;2�}κ�럷��$f6vt��]�S��b�Y����rw�S��D��9rڪ��帢qp��Cb��3�I�ڛ�4���ѯ7N��Q�כ�"Vj��D�%��}0�K)�S�P)�
X2���:��E  �d�^��J��B��%����d?��ew�U��V�d Q�odX�q9aNw�a��V��@H�0w��%*grB�:�&�<|����L����ެd���ٵe���w��5ly�ð�a!#��wBI2���>�����ҧ�;�٪3�9��A��C�{D�S�s��O:/�<Jq�1�e�)% ���x%nr��n+�FuJ����=�}��ܓ��T�u�,.z�tߊ!fV�ʹLk�q���x�
��y�����-����T��]���B����OQ(�uū�#y��U���s@��Z�Q���/J�3�p�YWv'�
����aw��
�P��d��(�9D�=>��b��(�$�..a]�#E���3^�����sV�+�ĩ9�U2AGN�����)�$J8�T��N9���>�H`��v�ȏ�=�A�:.��aT�M�J�=~a��ŀ"��������88X�PI8F��������q%״:h:��� ;�p�����
�����$S?�" �=o�u��Ē��q2N���e�K�~37�# {fzUzgk*ݵn���^ˈo�]�IO�TJz]�%Gl.2Z��L�vϞ�R*�[L� �ߣ����xO�xk�+��.��.�#��Eǀ�o��c�.g�#"Z�c07M��v�;(�w��n۳��F��ȍ;�� �'�{S��&�9�C�;�/���i�A��vg���d�o4��|@�eȢ�������2�k�F���0��dE2�\��E߷ViS�����S�b�b�E�@��U�%�h��$�t�6Q�~�Ov6õ�d�
W�2j�ީ��ƶ�q��.�@l��,�g_F��o��J#�j?����=[tX�<?��tL�-�l��Z��n��?����/�͊`��ȼ�ީ�8כ���1�Z� �9�� �- �|&;Q� ���E��,	�O�)X���� �j@%G�� ��녩���A��7�4��԰���0˷���R�I�r^�9��PslE.��f;vM�{s*��qI6�H�.ʶmFN��E*���\�I�V��$5�\{�;�G��)2�\:"� ^Ӫ;K���Xéٔ�,-&���!a�'�Q���5QR=�T?4Q�RM�x�4�ɲQǧ��}4��dD\o��iN��Z�E^_�c
Q�6Ʀ�z�y.�����jNDo�0H���&�hU-���n��W@5N�f4�Ū��"�w}�@�&����ۉ�)*@Fߎ��>�=@ĕ~��L��0͕�H�T��3̦؈���:pOz����������!�u�B>������t.a�?d"�V�(u�:'e���P(�0S�
j���!l"�_dN�X\~���(࠲Y�5�h{��_�R2�E*,B���Y�>���pz�H���M
��g���M�߆%[}�܅$�%l�vXR׫Ft��G����^v �Śy���K�Ɏ�V҉��l3F�ױr[ZQ��ø���}��r�D����d�O�������k6P�3�A�[ۦZ�������?o<��֧ެLujRt�	��&��M�K��M��j�t�f)��:d��<��c
;���6�A�-i�)�s�($�v�������Js�� �K9�H��>ͫ�U�GG�aR�GK%j��heON'�V�����Oha�\�1p"�o��
�<5�̓�$���,F�-�W�I`��Q��$M���xSй�_~tp`��O�N���B/��CۛZ><*���[��~��o�,��QE�ϸL
���!_��f�w���Izj��]��m@�_q�x~&���PC#W�g�Sk2��{r���!d��H]"0��v��o#�?���-y�w�p)�[sO��[>?U��a�(
V�gK��F´��U�w�v�k��<e��ﺶL�Hq�}�a�${�'?��\��Ƙcel�e/�*\t-@rxw�g�kO��VT~z�CݠkV4d2i;��Y4�=U�J
�~o&6y1W$�[�j����7	3�O��-��x� �!���AYA����)��H�L̆�ۦs��'F��a�Jdx
�ż�,=S��|r�_��zm ]p?���+aO�]X� a��� �@_.�S����W�����.0� ����]9%���I���n� ��w2\0����V:-^����3�j��a��3u}���@��4���}[����(���c�`�j ����<be����?RnCF�8���F�h���C��߸ �X�w��=v��	�?A��5�j�M-(���5V\���;ݮ���=n��X%c+#Y{)�� h��܆�FטΖ��=��+�	�7�D��I��O�]C���l��A
^�7���h�@p�ݠ��4]��VAa�q��4*�|� ͔��XiF"��9j��	������To-}�����!" �9�?/Z�7}F="�[��8�఩�=�����.� T�*6��G��rL�;��|���ʲk�0�Y�sQ �ߏ�'��]y)�����|�aِ>`O�LeV/ͩ;��N��U��Ae�����x���ڝ�q�_�!��cS�(E���#��W�mF9Y�Gq@�Eα��$�E9]���7�T�a!-+��&����ևY�߶�=����]�Uq�y԰���g�sGM�w�O��Lp|�d��V�����n��e/ �pP�ZS��z���a�W����uH� pX��V�؍���g��!���4��U�W?uaW���֟z�+�2
��ɭ��M������,l�;�l��Qz�o�����M�Bٵ}����u;\N82��3��0�M����4�����^a��<���BH0!�T-	i�77���/ȫB����D��Dt����F��JN�2o�?��~�v�
����<<�������1����A}(%�=pڤ�x���S<HN��f�;>ކ��HH!)Qd��%͆L)O؎q���u��9�Lw��4��tf2	�E&�d��d�t�B�p ��ޓ�/e�E>X:�j�A����~[MV@�rd-��{N\�\mr�����<TX�v_׆���[�vțT�֐'��Ŵ7d*���S(��N�`���:q���E[Qj>��	��xo���x�'c����gv����ջV�ۅ��#��O�8I�/��%p�-�J ΕmI��
Y/�Q����H-�P(�9O���J&2� ���7�X"�B	�����=(N׈�y^q�a�1�	PZo[gլ���kn��������^�B����\�1M�Z	촻���Y���?# �[U��9���|��!�R�� ��
�Ք-��KF�{���z`�:L6�Uc��4�h���V�)D���$on ����0&�d��f�<��'���\����eO�YM�&-�J��(쨀��Ɔ]F�Y_p\B�3��r&���d�5���k��q#�R�)cOI�9���[j�	x��/��t�����b�Ɵ�bM�Md�`7|��Ԉe�ǫ�e�U���:��=)�fՎl�L�_�C�T�tQ[��E�	���,l�腝������Y�����;Nc���ĥ����M��-���bئ9�ÿ��G�1N��؝���k�w�K��,�� ��_����Z3u�n�4���m%�o�*�����BG!郩a����u��y�����i�w�%���"X��ԍJ��5��(���1ݚo�#~	/��y2��%�r �\���� g��hB���S��s�qhe9sK_<z�c�8�\��cZ̒��g>�g�+Op^��\F$@��W"�3�.�� ��D��h��u9�����"�WW���}��e�B�rc�d0���
��/kʣ�l�	��ʅhx��~���8�%P�U'���5�i�y2!��9�=B0+n�=�'��?j���*�������{<}zme�{���+�Z��\���c���y���L4�ϙ�S�O��>����(��~Tg3��h��2�be���_��^��C��/K��7կS��Wm��cGS���ux��E8Tq�6؏�զf�_ss��-�>���āk��T8/,d�N��p��gL!�a�S6�o��{�x:��T���U!�n�-�(u}Wn�5����(�!+)�<��?��jj�m(댂�c��il2���6�E�N���.���W5K��.�HB��s�>Kn���Q��"��.�-ah��T�}�4bC�y����%h���p��4q�Q�xmF㜪��{�n�:�D��������Y](%Y���1�kB�9�Pr�G��)S����#��WQ���`��t��,�63��	�ևKF1~�?�r>X�]�IY�oom�:��G���s�2s9W�eBֈ�T�.A�����G�`[�iR�S�RpI���-�����\�mA+-�U�&T�K�����3%��ʬ�0$��q�*d�l<��k)�cN�Pپ	I]1a@:}�-.�hk0T��*�O��	U4��2%�A��9���D�ީ�5��3u:"25�$Upb³��tW����TO�b�3�-)��̉A�Z����k��k��o�o+�~~��"y��xk�����H���NFwH�#.ݨg�P��Q.\	�/;�&�U)��-Hz ��%PH��P�}��U���I*c��{��t��)�,�P����]<#Ĥj�Q�k��Q"	=���M�ŻX��%�+�p��-!�ý�����?�^��X��Ylf�h�O��s)$e�9u,�m�MJ\�x02�"���q�2�Ѥsı9���Z@��5�^_�M$4����K;G�|��E���<�.�D�v
��	�t�X8�ǄƋ|�l�⯊���]YU-��oVU��(�7U-F`��ۮa\����;�I�:���{
T����g��|$H��Q�mi97-!1�mW$N"�"����z���=��b>�����Z�s�L&�ws
��'~`�w��@!m
�^1�~�6��7��ܵ��C��k��L�g�B�ĺ>�3��Dp�v�1w�z�H0��S�(Z��ŧ3�8�-�4�f�����	%1��M!T����c��n���qcak(EVZ���<����i^�H"�˂�(/����\0Md���=ݪ~Cx�0�&��ޙg����J#3H��=�㭩�����')��0(w�B�/�����T�Ps]a\���	Ƭq8Nּ�P��c02 �-���HY��D=�t!��ʅ�7���2���h�r�}i�U1F�·ʇ���nJK����;8�]��a3\>O��h����ߋ��ԦIN��:�tJ�����@�:d���/���f1@��	r�F��z�zqdV�d�azc�zL�JZȢkJ%�^�܂357!�+��;2��32�����D꿕��*�A��(��&�]7x{��3ڛ��D/�yq	�Lp}%b�c2,��)*�m������;y��n��s~+����ͮ��PVAV���!q�����_@@OE��DS�:fXuBj�xG����CT�gηn��z�zD$�@�Q�e$�Ƀ�:e�3�X[�n�_�E��o�3t�W=]ӄ���@JiU̐�%�=�\�{���7��g�-6k��$1#�V�ٿ�����$)~U���&�n�0��I�+����]])��(:��tf*H�:{��7*�X��[
�8�d|7P�����E!���=���MC����=�Nz|�,Sa7��uk���E~��\-�8�.��򛨴n��D�`���t��fX��6������[�!t�d���0)�Q���2e}S�������^Y�!���q�-Qԭ�ED�L�<]xߔ�Tj;��/b�ߦ���L��<%����*���Q�� �C�j�į��ܷ�-����������%��}O*�&A,��=�C���U|Oh��'�㽞���&�x��l�𐇛 .�?�P�y�0�q���늆r@�>��	���ϕ�ۚ�o|����:��MhV��d {Y�.?�$8>ȀCk�����z�o?1�#�~���N�I��a�a9ס��{�D_�7"�S�=��rK�m����8ݩ7'3Cշ�a����i_�Wם�����bI@JVc(?���i�@����6�u���G4@�A��q��3}�� 饽æf3>u�r�|������.͵�W'���JJ����^
gX�&a(��� ��[�؎-,;�v��5��ž��3F�)!$��N��n{���^>�*�3����P���3gM��p�3	����Y�M*�#.����z�jdQ�hbs���<��>A�x�d�`����FP���\�]D��Y_%��
�����[z��l��?��*�+�;����7�[I-�t�}�K$Jjk�y�rr��N���m��⤼a������eq�v�b�\*������{!	��GY�4�6�>�<L��M�K�6���F[��-y��(p�����ՙd�Σ�2�O�45/�Q������6cc�k��Oʩǎ 6�K?�&�:�p��B|�?��㕘������qh3��o��}$t&C���e�٤-���N�eHY1��͵�4���g����P*�e93a�rT�ԬJn����TL�ǀ��}3��Z�:��C횑�S�gi!�n5A��z/d�b����r��'	��8en��ܺfaj��v�
@�4�H�{��r��۶��J{��Z_�������h���[�l0o6��K n�dn�'݁�����/@�(��-�s���_�B���Z`���g��8;ȗ]��bᓊ����8��8
�� ��#�ѣwk�LYEdZ~��e0.sX���S��WB�
������ʙŘ�K"r�@s����oa2dW?��&��Bs�a��O�Vu��vU.c��Պ��r�."�,_&�V�:d:�.&�������(8�ʤSl�s6�f($u���vn��5���Zqmv�o+4?�����kRSt��I9�^ƵA	5i�w��}\0$h��6R�1������q:�9�]�2y��~��}��(k	��~�PB�ħ�N+j�!�+?iz�Y�>�����|��6�D�t�B�`�i��cM��b}��<�	�Z���b��BA�$�~��PN��ʄ��z�)n/b����L�kB;ṋb�7ոۏ�H�+us���&�����h�G5��uO��g���!���I�)���M��@~4(W�5ۗ���z�`+F��&��8��	�RW�������]K�Zl_Q"�Z$_�v~
���B��W\V��5�w�>��U̑���/�3Ќӣ	���@�mq��'~B�\:"X*Y���AUZ��'}1������6H�r�(��R��_��_`��'���$j�>�B^p����ڽI���T<驆x6a+�q�'�w���z�h��ǱU(�HG2(Ok�4�oK��*Y�}A�e�K�Ǘ�8̒��X���P�)�1�v7�q�ק��6��,�^��|~��!�C!5
�x��Ҩ��h��k���Ӂ>{���>WQ���=���~h��x��A%8�F(�w�hڜp+#�hU\>�K(,N�۪%�����c�簻B;��tz옶�ٞ��/ �$p��S$�0�N�y�G��+"�'<��Ȑ�R�?K��y�w�޵E��yY��w�ݮ�eĨ'W��z����d)�aC��F�� � ����kac�J�ڙVd}�yX��t%?&�y|��.Ɠߛf��J®�����K���;,�Ǫ�w�*������"�����Q�W�k>�0�S��S����Pf��%���<�8�$���F�R(�=:��"��ʨ���t��@��v��k�t��(�mo�ZA��6a^��F��z�r��񇉹�!?�X�+�m���W����·�HD�Ç��d�*���1W��_�XӔeO��e�i�Y� ��A�p$��}�{e�M�>�E;!�4x�Ś��+���d{j��'{�#S�zL�6`c�^��p�i��q��U�M9�;�*�uu��HzC g�.h� h-n��Nx����O Ip�m�*���껖�n�p���� ��BY��=Y � �b�)��O��^�ש��%���$���萰��ɵ-��q꫉�;}Q\9a0��gjU�)8vkH��{��:mt��֨]���yo�@�6�zj�o͞�ȷh�(�~E�K�T�6�x[{��d?��~�TEk+�<�u�;pD	#�M�pvFDB��u�	$��ΤvKfٟ4���fa�XBT=��և$LZ)�h�l���j�oO�$
(9C8H'G�'SSGX̷8��.h6�w^�-\�G���6
�QE�YGS�_�>g�;��`t;9%+4�~GϚb1�,7�~R�@�{�]J@Ux��`+ֽ��̾�s�,��؈�*�癋y���Q�˒��т�D�˽�5��ۡ�iH�-���C��Yں�
����)��,����d�%r�.�D!���'	?�c�D汬5`��8ײ�e(���5A�5~��6��(�������U'�jd\�rhl�{\�ӑ��y`�lB�S��Z�biR�s���Btk�&/��%h�����Z�b�QuoP�_ *��*�E�S�a�$�F��G �բS��J��q��Q�6�O5�{�@�6���*�B/�{�3a����kPvP|��M�����# '�
�!�8���q�N�*d���z���ls�8I��%�kgy%<]�Zx��4w!�8W��CQi��rc�2�*]�Sf���`N���ΔLo�Em����{<�y��s�|n��Z���|c�[˛����l%��U���q8*��N�
,Բ�9W����K�{��������^�=�(=l#m<v��Gz�Zo�l����f��!���C�2cN���1�y�3���+w��'R�ݠ�%����T�N:�M�	�w���.����B���!�\�lk<�˼x�*G@v�C��ҟ=%^��j��L,���f,��"i?F�Y�:(Ib�Q�%Zo�{N��%]��a��	�� �����>J�@�l"��_�JV�!d���}:A���cX6�X�*�E΄J�LP��9_0�*�T� APNV��`�"w��Pr)Ԑ�`�z�A CKn����3j63,��n���ܫ�����6��E�20ܵ@�6�[��	X>YY��#���B2�R�����ݱ1"��c+N�;3B�H$G|����n���B�,��4�L3���t�5�Y�~�]zÐ��X:���k`l��gy���e�x���㋧�xA�T8�}À��m����~Y�8�9y��:b2_�[D9��ގ/B�Fװ����ΤB<�t�R�Hm����.*w�S!�A��2�~���c!:#�s�-B��(S^NuF�����Js�~�%Ѧ��B��yp�<J�	�� Q��)�L`Yf�.j-�GG�<����-K��`Aił��6�xe��/��&;���huS�m)J8��xΰ��_����+�T�a=D�6�&�"�	:���yy郆����T�����Q�����B����G��uO��*"�E���S��,�!�* ��0��k�����{�hM&_Ƙ�B�Lk�Y'��#�Ի�&8%��>��Ӷp�c�%Y6�R���5�KPsA	��f�eٻuf�В�DH��b� 'ꛠ�1�����넩�G��#�2�t�7>{iӝ�57-l��b�h%�����Gy��	� ��Ǣ^g, �*��>A���������-�x�6y�M�-�B��F�\�=^���l�s(X��}�CSz�\���4���fl�XIw�����u!���ڧ��{,۬�L*��~V�&햰J�����M�RI��#��7�ruhY���#�̟[�PB�D+Y�+�-���j�Zą���dQ)��|����~�H$f1�S�|I$a��l3�De��:O�ճb���77��؁�{���&FBNFdE�"/�?�OZTyp.�����5�,'%��:IX]+H�W��oV��$<#\J�`�mU�d�-���H�B�gb;c��k���%��]�D�zV�b5C��e�ˬa)6pP)D�\�!��y0�\�����"���B+&�W��9׏��d�~�l�%M��`��ld�(����Se`V�Gg:���fRWkAӁϔ���u�
�HbI0#����8g��ɹ��(sV �m�*D�+�M"r�L�H�ZBo���� �_q��RߘoFjpt���A�$M�l��|q�4�+&�f���
@v&s wXF4SB�,�D&+ -e���'��TD�	��S)���U�l�e�� �����[��1T|5ؾ�Qoӂ�K��c8-�|l��)���@56A��i�4�� ���b��U�vh'a�p�`*\���a>c�U�'�;+�����Pm��zh^a���ɣe5���$Z��/F��I"�dJ�:E|إ&��?Cr��Qp�	����7�j��SS�|�5�=���΃�э�|��+�E��y�v��+���ݪ%��J�I�0t~&�&�pb����P���ɍy}���l1�d����!c��Ԯ�qƏ���S�44�֚Lm��J����D��{���R�k���U猌k𕡳a�!aL.�Qh�<�<��	�z��|x��X�C��:�2ޱJ��i��d������?~C�2�+E�|���П]4�� Ҙ�E���DX�,��ASh�^��0��S�3��5m %��Q����/����|}�F���:i�uj������Q������;�D��&f�/���;���xNbR��*��)���W!�C�n�>Wo��e���W)�F�K,ZV���i`��=��w�[A��U1)̊S3���?�����	x�M�C��ھā${F�C)s3�� ���1��Fa����.�;�׵bϕ���� 
�ݽ!T/��!d�8�w,L�SB���X�1�Qث���j���2!����Ц�I@�$�8e�4��q p�T�.B����h����@��Eܮe��D��p6�Q����%�kw�j�P����r����Gv�H�硸�YD�g�i��>ː4LI�]�o�q��![�8��z��2�{�w(������%՗UG���=}I�ͷ&LD�(�;J�r�p�����)�
ąI��kI��������łM�����J�=Q]�J����t�m4ˑ�>������s*�J�ud�Z��0F��r�}I�ۂ��M��e	���:�H6ͥɲ#��f����dP�����-w!^a����s����/���@�%��$6P�T�yt��/_���4
��6������oV�F #�Gc����0u�������]{G�'R`T���4�0aj�Nx[@��ה;��ÇG0G!��XE�$D����fYA�y����O���V.|�4�����+�#	E��F�خ��5���ۨ��� �:c-�{�@��ϵ���$!�c��cDߢY����+P-&��rF�i�T� ��^h/g�e��`����k���u����OJ̃�'��eHm&����[�N�6�=���ke�auq���Մ��6D�{II�X�v �+���j��p3�Yٹ���oOW����\l���o5՝��j�o� ������rOc�h����XA��}�,|��i�$B ��G�gYd�ĵ�Ia<�������l{��2����VQ�6��4�PM�2���0#k��fF��#ͅ��#��E�(��T��.��8߽��+������NK��|90-ɽi6�
i���7��1چ�l�� X��V�,m���QG.�t漏����S��<���>B�l��.w9��!d��m&�y:
�{��s]d���P	����NJ�G���Ԅ��=?��$�;�#��D0rS���-sI���`��EMFb��p���f��X�b@��E�HT0��L'��0���s��/U�,�G�������a�3Q3a�� ��H�dJzf^��5Zf�'d�ne���Z��P��s�H�Z�!��SY�����A�X]5���z͛�K��/]^E��M�uc=�VGO�� ��%�[�z�V(3�{ �'�)Y(_?�u-���*�^*ƚ���v�VL��z�kG)֊�Юcw��� �S
��)8��Ԏ�Sf|�(�����R�Fl���#_�.�J���lh{�LE��ȣ�.+5^E��,��7{�s�)s������^��Z;&Z�Yj�F��}�1L22���oEz��rCE�6�k'۳�3���C	Rzt��!Ja�g�4&u�L���ӻd	f!�ln�)�
Լ��U�V���K}����Z0�ì�d~e��'y�d������~P��_l6|�xg��Si���#��(߫z�7�X �Q֥��Wa!����Pa;��R��׃wa�EEBbX>��A�[xEE����*)ͱ�*�´�W#,  ܈l������U<�k��֐�ݥ�e��y�sI���ݷ���s#����O[BB�/�X���^C���f���JĮ�Ov���Q��ۀ���%_��7a��D������ɼs�5/����Ui$��^��V;�	|�����t҄�!ӿ��Ƴ�ˊe>$�������D���D��=�9�ؗ�q�	�os7yr�~��F�� �I��>��q\%t"<^��2M�ߨ���L���8gqŏ �kz�]��R��c��7��ڤj��'-��w�`ș����u�D�!`,���v���2Z5IGŸmćŔ|�9%kT͹���A]xN�G7����gb�F�P�uhͨdC�`P��H����=�#�X����,�e�D]�!xF�O��&�%���6���n2N��2�FX� R (���c�ݺ(KGz:BZ=�����~Gs�z���'�*���!;������
���B���Y��4a&�uZ�7ŋ��`���<G��HQ!˭_��w�N?]A�U5�M����sR� �7�v7/g�l�aŀa
��F�[��	q�`+���CS�a5z�{P�#Q��ca8t��bF�m��S]V���k�b��sEǶ�Cѭb����7�wC��	����#n8zm�|����r��a�������������Q�B}H7.Ɵz4t4�Xё<Q��[(ǎ�����^ �J�ʙ�rt��-X�(+D`�j���9�'�<�q�92:�5�r�t��� ��E�<��e�L�f�svB�`6��0�`�s�p5�h
���t.�Q���+T�e|Q�!(�4��I��@m����C3���@s�6��i��<���qd��z�	L��X��؅���z��gۆ-���3��sqP�(M,vd3U��Wub	Q�'ɱ�a���}Ժ��PD�E��xV3&#
�j��{�h�ĭ�ӏ5�ޠ<���ˤ-P��m�P�.��<*�6�O)��Q=�%d_��䳚��M��Όc>��.�N^w	�����Ri��i��h����T-���%qՍ���TS�%\fq�|�n���u�Yߦ��k�~��6}��$GK��AH	�ܲٝ��6���ɟ�=^AD���g3��{�L3ճ�'�� I��"�f�>�g�%�o����i���5ܫ��"�o������5���sUS�qF��JL?�������B�LSʋ�g�7V�� �ľR�0�6�k����q�m���}�l�+g�l�Z��#`��4�S��ܐ']~K��
L�N}��/�6o��~rt=���|��p(rtw�zaC�F�s�o'�K�l��������sǢU�'��"X�X��n�&�>d�/��j�0X�Y���$l�U�V�B����XW$�N��S4����C��Ee��,,�e����B�-�g���إ�����wR�U��N[{���}��*����Ą��F'�/Zӓ���������
�K[�Jj���y"m�	�P:�%c03x�>=N���P3ʡM�^Ճy�^du�7�j?��1�E}U�
��+1��ݵ�CO2�-.���u�\M���0ƕ7�'�Y�\,�ϰ��b5����~·�G��tI�=�9�4��x]ѕ�������j[D��/1�}H<,��QOZr��EņS����k-��=�r�\G�	G�͏��u�BUT�"�����c1.}�*�,vk �#�l��~+��k����l�/�L�x�-2�ſ�p��YD�P͡T�f��J��������������۩٦q�O��c�8��ɣoY��;��
ξ�͏tɏ�i�)ּN�L-�2�:ӝ�Ɖ/�YqOKSI�p��y�p�ެ����9��6�܂���
��������)f�b�w�Yz�?���C�]����D���6��~����as���O,)�
SF��M�B�u78����� ��;%� �AWhjsL�NO>x
ۄū��.1�on�2����mD�f�=���"ư�ix�9d��L̰
5B���IM�t>�8�ɲը�7�G��Ctarhe�?q�.���x��l�����#P�6�^q�P;diĥ�揸�c%L�سA�h�'�j���Y�y�-�����K�ń�f�2��^��	<�İ�a��ƭA�"D↌,�_l�qJ�<��?R5Jq����r�{7�k�K��Ǹ�{�w\� JkFOc�I��yz4�5�˨��ZF�z9S�k�4�l���x�X��k��҂�ҢFy�x|�+��d�H��k򩐠�Tb�
�Pt=5xBLd�S�$,�Q���,����k�Q�!��H��1�B9ZVP���[�㶤��Q
9�����P���<`�/�i9 �� W�z�w�=��B �1����:}t����O�Bs�� �'ڬ�؛`�e� ?T�,�:�hLe�T���7>69�~mHT5���)1S�����	��b�0t��۠���4�>yO�_US��օSϨO^��9)���ĒCTE5/Yz+�n-zD��T�`��aE�ׂ~����6#�Z�u�NA�㩛^t��fR�q������iI8�sR�vQS$� 4�}P�w�|6C�R�[Ʃ��*I�"R3[�^]�`���S0 �VxY`��Cڛ�2��f`f/��5(M�ץ�*`L�C�	��B;ܘ�ʏ+��3ů��u}�Қ�%��@�˘[����&�ľ.�+Oo��Yk���a%V[����y���g?R�/F���Ge�7Ic�N	�/C���G�[�yP��{V�ߙr���N��<2��&,f5��2��AF	�9�..���Aǰ6�2�㿐6�jܱ(=8C�0���b��{ɒ?:���;��u��|c(*i���E�N��i�+�G��,��\�]m#*�FbC��4��-5���(D����GP����2t(�f��d�����B�]�[�d�{�q��Y{��ئj5�&�^����_�l�AC�+���;�,���8.4�N��s֤��l�h#B�uN���� �=�N���,"H��I�/b7��3"����� ����W����?su��}q٠+,k�]p��;u�p�1����jvI��/���d3]�	'�a���Fj�����o�J���X���*�~�\wl���o��L����=cr��zv;���`��q��~.�w!;r��ݢ�きn6,|n����(=:A$�
������騐�b����(M�
�jn��e)gE�)��ԃ�</��Bw�bQ�o!����1Ѿ��@����N%z��z�?�kB�����
Q~�JfF+t*�G������O�{Φ�ER�� �G :���yg.K[Xh��V@ ��
��~�"�D�i�Yb}v������̔/�^xy�+Ɉ)�^Qfc�hG����jV�(��Qa	*dߕ�^�SܝM���5?�!��#B��0}7 �R�4�؂y9A�HV
ch}z�e����8]5�yPSő�⽵���k'e�fGa������t�2p�Z$�R���b9�:'�n-5��m%����oj6��O�#�a�
��p���
m�5��Rn/Cm2+,5�r�gP��g��|�Ƽ�ɥ~�m�����V�J��x�>�oa�"��|��v��M���#��=j�,����?���h���iH�Cn|N�D�`+c�A���L����836]nf
Vb��ׂf.��IR��7J?�b�����k�aYe��ɨ�_æ-�H�� /�2Hd��fBp�"��P����Џ,�BKH��Mu^R����>�3+q�`c��y2���uŋ-�^B�~y~�����5#Լ�^�yR7�k���_�؀ ����7�#b+�wu��1j�<�7��9ܯ�_bS�r����R]�6�֟��:�>�R.���3ߐ��]�Qcz��n�j�B�X��3$�V��C�d4_��mĹ��t���X�A	�p��a@�ur,�44�x@�����XmwТ'��%H���O���r:S�-o:��i@BF���Kӻ��Á�PZD�b	��<�p{���$��0��`4)���6�E����	���Q�'f��4��Jλy���FN0�V��،&�OO�[Z)��v	G@6�#��z��b�����KF�zt�*����	�rTӴ��(�42=\��ц��B[�u���o���g3����<4$�D�t��vi ���2%\��:�A'B�'=�.����Z�`��b�@�W(�Z�UR��� ��q��eq�yoɗ���j.f���~�7�h�A���A�$g�Vs7�/��9�;1ц�PRw��q��$9.�І����S�h�2�E�����O7S���82�é��]�Dj�oa��Z
է�r�T����V���������X��DfT;z)���'B�6���O�2�:��Cf�J ߇S���O�g���.�-<R�0� ���5��.���XY��l�|�_p��(����a��|QH�8K�>�'JK�@�GL�S�ggbPj����0|� |K"�
:�<�W�RC�:� ��U\��2�3a
X�#��k<[ɮʆ��]0��x i�p�c��Nt�hӼ}!c�T����k����w/=x$0̉Ƚ��b��ۮ�62�=�f"��`�7,C���7��"8ދH�ABq�i(b`y�;Il��L-��|���[l�!��=k��~�2�]���I����,�,��u3�3#�]+O=�}���� ��^�S]���:bi���!�[�5��W������Y�#si����D���8�#���s���~��T��*O|f,��'x�ȭ�-66{2�8��h^�(ʒGU`a�(rrӑlFz�
ܕ�cK��uH�>�[�Z��ǕtP��m���y�:�b�oOۊ2Tz�`�S%�G"n�t�x�&�Ε� �� S��{A���ŵ,z�(���P���L@,g�k#/]6�!f'��i�ȃ��# g"�/X��oR!�y�N�Oc�ԖM�%-?��=ce�T ]2�ea�8�����({�[P����Nl|�g�Y���J��Y��,�oռ?VnȐ��mZm�
v����Z-y�:����Oˎi[y�|����jb��Z�LW-R��������A���(��'��R5*��tnK\��~��"].�(ҊU��6@�}��8;P"a ��+��5��r�`�`�27���I��W��Sr��|bV\1;�D��;Zp�T�Щ���Lߟ"<蛰Vu,��2
�,�$�I3��J֚�~
����_3�[�a
㈕��u�:f���7��n�Lu�xs�&�a���/���"��L4d7��;���Z`�sh��"�S~����j�*�:���.�d��8�?��N<����K! �+?s�ӧ�#Ȫ0��AD�{8�U�.�$d���ٲWB�p׫nV�B��~%Jǋ�6��*�<���Kt�����R�Z��	T;k�:6���4���
�ES�_���j��\Q�]f��v~K<�x�=}��hM/Ġ��L�x����bc ,,�y���.��ܑʰ	|�c���\�ۖv���$�K����v�5�:����f;f���]άTM����	ه��z޸�7����|�-K��`?"�-����
���mm@U����/jPS�����KX�Ԍ��Y�$3kq �Ӟ�1Z�j��P��D�d����b�S[��ڣc���T�)K�F4D!,�4P��8XD2u!�h�.99!��mR�m6���ժp4z����[.u� �}4>7���>�9�s<:$Ww����Y&Z%e@�f�ǚPc��>�G�տ���z�f����e߶�%'�O��K�z9D���&��W��n���Q_��Wa�m&r��*?F�� �:'�A�`q�b\�ܐ�SHۣ��d>A�dD[e	�g� [dP�M/ϟ]���4�����Q�6��<�>5�J}~2䭇���XߜT�9���y�����m�BC���\����}��+������ �n4)�q�p�3�����%�4�N�/�ɫ�w�s�7Gu�� ?�ݼr�ۊ��m�=��
!�%ȷ�e��!��h��Sd���(����{Mæ�=�=͐b��.@�~9 <C�zFU���Rt���5�����3��S���ɠR�Fx=Lw�`v��3ƺ����*����[�^�\(�ӫ%�f`AD���3|д�L���� ��QV_N_��\y���T�Z�}\d�����,9a�+P�ج�I�aאt���A�]rA�ݐ	ߌ.�O��p��i�zKc�eBu�	;�'���\!�j2��o��1��lbL����4�¤_�'��f��7ny�h\'=���B��A.�A�	2�֏��(f�јwɶj��&�v��ꀆ�s�l:���S�LG�Jùfe�z�X��%�C������$�2	&_QE�	����FC���|�c3��.<��wZ���iO�s���V�f��e��Ԏ�m%�� ~�x�c@|\��s��C�G>��N.�C �PW5p$q9��u�>/�VBF�Q�Z���*�]��,P�
�U�O�>��Ud�n01�š���<��Q ��GJ~-�МҐ�ܢPK���;Q�z��Vxce%Y$��o��|1����@������
2��|�8.�l��'�	K�A��X��J�s��+E�����r8���ۨ�\&sI)nfT�Kt��>��N��;�h��j�,���o"��]cf�einYx����B��^%��T
f�1|ub�x=� 	��>.��rX��T"F�7C���M��y9� Pv#4&��G�Jh�a/�{�_�mt���T%��c��uȚN�ߋ<r�XJ�R;)����=r������FJ}���������Dz�$*�:S%$�N7������pu���t�$�����[��
':����I*��C�m@�tq�*�N�қ�+�5����l ��J�t� ֲ8�3�V��z�V��{�O\�4P6�u��D\�\RvkA��q��S5`8��f ���޷��V��5܊�.*�1zJ���7�JL [�	�u^��9p
k�~�E��?�\����!���Jҍ��nk�K���R����G�²xN�.�f��t�����o���ϋJ G�����M�W�,7�7ۮ��5�<�^��4�kon�m�t�6!L�XҶ�4����0��Y�0��N�[<@��%���LVh��-E�WG�柳�����se`��[���˙�d5��WD`Y���?P�A�FU�4��y�%楝����	A����x�y�U\�9�q��
����n����q�v4I�j6X7M�O�����|�=9,\��=��VFU(�z�� �m��qp��A��%���q=���f�1q4����q��|#ס� C��>�	_n}\�\#lP�ޥ�m���F0f��Ď3�ng
�K��#x�n2�L��b��ż�NZ��͜ʢՄ�Q�{�7R�XK(}�펉���Oa.Y�I�y�s=�k�ۡ���W�jѵ�t~�����g{�K_
=T7x�T�o��.��`Ҽ�!�h�Ij��f������H6�+[�Z���8ɓ?#Ȓ�f�!3u�]�8s��J��HA�z��=�Ǻ2L3��	���_e���"V�q�TZۯv�7�J�I�!w��P�8�x��?<�IŸ�o�x���S���l�J/��6rn�7$V-�K���t�*�9
K9�L��B���݁�&�+�..�t�V�U1Q,�2��	˺�z�l���p
�7n�4؊_;�=�4�5 �ǿQ(�H4I�A(�8�ol��.޺t�u+������%�E7N���a���h���DN�+���z&����@h�3� �s�S QH+^�dGMˠ�9N��V�#$#o{�z�j�&���|!��0h�L�^���7���,�qpD���Daml�p-`{�N(׍�]�X܋���+�ev�^��2��f��gzzx8UC�>��
$Ɯ��f���խ�(��|�@(�ݕ���5@�{���-Kf�)���-�$��(��D2�8���d͊ ���-[?M�:���բd2}͝�|�GCLc�m����.�Ҡ���c&CL
,̢	�~ ���8x����ez��nH���|:HFV*�P6�®2|��j���>h?n]�f�w��9���J�ԓ)َ����@���=�̶���TC�{�Yz ��ۃ��K���#�~l1��j�q����*Am�)�r �W�����/eEi����S�����+m�!�U��в#���Z���xy5���o����� �z���^��������=�w�26����S�uڿ��_�6��)��
��ǔ���ϫ;A��@̆�#�﶑BY��jk~��A�E��%s��U�!��x��b�@Y��n
@?[������*�ۧV�n��(gW	�k�b�^�$�rh/�]L�V �������.L��g�w}tAR>�?�ZQ0O�����yG�t�e���F�8$���RL)˥����Z����-�����+��C޶]���%YZ�f�!�7��[Q�Xvrr��W�.q�Ұ��l�m�����xy�P��lbj��
X2(&�ƞ����*�x�oQ<�gx��Z����st�
�]z���!2f�I��:Wa7�G�a㔊¦�H��W&RW�"�.<Tf�2�i�� |< ��7���q u�
g�	�����t3�s ,�����P��v�W�o���-J�`�6�T+S�e$a{� .�� ��E1a��-GB*��c���) -��ե�$j㵦Qq��� VJ$׉	�*�e�z,(x�n�\�k��ўAt5s&��!	<|N�]r�����lP>f+�E�`�4㿬��qaӌ*��@��u���75��l�ܪ:�1���xH�Z�J�	��	 ���R�%���*�db�T$���j-DEn�˚�Z��Q�,�h�Ž�|c���Y�L=�h�f��;񼰳����%�+6���r�i�#0$���aXFf?��ڱ'|m�fG�O# �6�$<�q?��{>�K�Q�0M�[�|wXZ�2;I�����ʛ�*m�ne�3?.=QYr3��dˡJ��!�ħ[i����u�e��9�j]�Pcq�
9������IM��vߎ��ܶ5Y�$R^�{���������KU�+�7RҤ������Ww����诤Pָ�`O����gH3���hb�,�dըhMc��L�o����/7L�GHsEȘ�[?�A��z�٩��V_
9j��*�!o>�%�K��*r�\{�!5�U|厌l��Q�v.xL�:9�O����&s�n���A8Ty�no��f�'�������b��u�@�DD�NI��̡�\���T����8a"����*Y-&�S�}�x�6��	uJ�Ы �����S?��P�`5y��C ���,np�oƨh@U�81�G����jw.�� ����E
�n�-��E-Зl��:��*�*��(2h%W��U�
�&���Vs+���w��13I�󢢚�w�L:��a�G�Ӷ�;�oEы芲��}G�6��U�Z�ui���ds�ά���̴�P���J��Y#Nݗ�c7W:}���*��Y��L�&J����F��7�G
�+SuNb�ǆ8!_6�>����y��1~G%�R�"Τ��$�w���I�M�ai�M�ܭ֘�����M<��b��vy÷��!��w���HY\Yy���U{��dm(���ɝ���^.���~P�D�S#���xl��@�쀧��E�>�h$�ˏ�nLQx&ɽe�U�K��H9ٹ,����e���c��?+u'��F�%��^W[Q�<f]�!r����>�w���,CP�>m��,N����T�S^x�'Yb!���������´�I������j��k��KH_|ܝ �浕zriѳ��i7��	ƈ�?S��
���-�ڷ��r��f\F��/�N���ŒB�8Kg/�$d����?]�m����Ng >>���+z���B��w����I�����Ju����Y�_>�+���O5��!��K��J����m��\�8���u�.��^ћCa�Ta3�S�P��sc�H7��<�0��L�)������`��*�Rp��n�mƘ����MLn�2��xū�����A.��O�4�u��\��n ���Y%<���������<q�n�y��HAǺ/;�� C�a�k**A�2d�
�H����D�yU	y=v��v�A]P!	LN=b�n"L��Zqv���A���2ʅ!)��*���9,#��d����̝�2�Q�l�cu��xP��"�nuM��(1'�	��Ԩg�eǮ�u�	:�f�b؎:�u��[ʪ�IC�2+�V�GM� ���#��B5L䐸����;��_��%�3�RW�ޖ��X ����M��:�	�`�/@����}U��E��0�(�����HtQ��������h�E�L���$�`�%��U�#*ֵo�eNn�&k>=����)G��x[�ۻcP�x�4�g�A2���
�D���lY�b`!���oxdgz��)�a�������G��n>�!-ri��I,3MøD�V�(�C^�Ռ��a��6�Ƭsz��D"��.̇$�[�˶%(��\�&�:b�Cٞ���^LO-��C|�+����Y Q�"�!�b��/I��QT�Y�<�{��`�`����Xw#JI=�D�����[~��^K\?��H����RU'�t�ǯߜ�u��kE����f�?7b������ui-l�p��Wu<#k��2��Ԯ��V��Q�GL3���o�{�^�#��81ܦK� S���ȞRt7�υr �
��}{Ǉ�.ܝ�{S�#��ٟ�c+%��lP1���,�x	d�ғƐ�+]�I�녋@H 3b@�M�玘a�P��d�㼺�-���>�VܺA3Ȉ�����6���t�'ك^V�����_���ơP0~b*�8���p¬WD���ȟ�1b�c��l^k&)��tLu&c!o������	sK��|�y�*�[����]Z�K"�7�q����L������C��4^�iĪȟ^Iur�1��#>SnP�_=OH�wt��yAGiOMt�k�t�5��M(R=�GLqh����
ؾ���}�v����
I��ܢ�'-hy T��I��TC)J���/�f�W��(���9m��Mp]�]��٦�DU�9N�hU��"$�o!�s��h�W-c?����~��^ĵ�����F�=��P�����)t	�ٛM���ςk�p�i�9@��E���l���>��p�����;�̓���v�u�2��~��46y\OGȳ6�ڶr��t�%��Z��kC.���1��� �ͬ�ۼh�wmĪ��k����۶4��ON��|��yrm�\Z�T-o5���S�v2��MŴ )`J�aD�w�����V����M�<�_u��x���bع�2�� �QK�f�ZI��,*+S���rЄ�>��������`����s����n/�+�%�j7�|��=�1�ؒ����ϸSM��̖.�W��v�-�Ph�A`��,#���q��:-�{@/|��i��ǋ��T��o�����;���~�䛢�+fv��Z����F���i�H�h������_�Oj�-\@૸�Oo��Gl6>04V�<��Q�x��" �\ �L�Y�٤�f��$�ēQhi ����rWB�i�9���&�߫�v�$M�QDE�a_a�PM�N�E�PWdv@�S�=kS�{d�0�0�QR�:<���&?�l����u���;F�-0�rN>~�x���V��)�f�K?�[��v��cwV�8�@(C}��FM�����/��@�d�E�ՑM̕4��K�t@5ty`>��G��I�M�����_§/+��Fw`��,X3&QͩKcWaq3����g��$B��Uq��f:���Y\z��w�{@���Ֆ��v	�A�