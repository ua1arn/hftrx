��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+�����b�k�t<n��!_^|�0C{����+�f(���͋{���'�*�
��(�C��5���P-E2"*��t�[���E���E��dZ��J�pfq����@\�m��_�(�#x-�=?뜿�X�(�N���J
�\;&�;2"�%�ZV��,�؞����g*7�����'l�������`h����Wr���!8�ROX�f7)�
� �OP��%`}��QB7��I�0�b��<���KdD�8��^�R}�/��"8��lo2���[���
[Z�%$�w ��ah��0N-23>�h2�i���[��ﰆk��me텦�<��w�f�'u6��`�,~5���8{?���jJ\���_x�pjsԎYa�4a�]�X��2�-*����n6�4���Tl�D��^[Q��I�v�/�v����xى�{_����A�GG�*
�|�%rL}����� �(|{�u��g5��&��,���AЫ��\�Z��~`�1��ά�a���,0���cD�3+���P�(X�F(�ܠ<.�Cy�x�L�q����)�~[b� C ��z�շC\��|� C3��z'ٿ�{���UȔ��	]$�qO{��Lù4s��Uȭ3<l~�%��ژ��0[0 ��^!�e0�z"���rq�zO�P0f�i��t��`d�ĺ�p�ƃFU����3�JA�NQ�=�)�c��,��z�H�y��Bl��Ǩwi�[)U7��C?o4|m³�/�k�-�X����W�J���#_(x����p������	�c]ԞM��oA7!��RkJ��WX�#�^�]}�a,2��f���K �~���HMY�W����7�e?�/���I���1k��X1�i����R��N~x��Ջ
����<����$���*
�o�����t!��s���N.`wd\ n�h^Aڼ���9nI�xLO��fU� 36�5���
	��������OvE\�!c#�� ���:��0dYֲj�w�5��./�Ad苪L!�S�ݯ<�|Q��d�=�7}>�[����5$���A ����KH���}6��i���y��]���709B)�f�����kl:G+mv�F�������28�O1@ZH����u%덳 �J{-��@�����*c:%�V�~��79����� �v���{~�����)R��5+7�U�ޕ�eJ��|���67F ��s�b/n{�2�x\�ʡÀ�)hmN
,]	���q�Fn.#`O*m���8�=]��9� W`-+��ʔf�9��ߒ<���F�I���H�����.���ױ�Cp0��X������#������|�C��:>��9��̺��S��.<�,���K���*a!�u޷��9�O���M�*��Z�
 ��.�U+�K#����rõ5�=�1�>�x�&�a�-��|"��X�4���ue:�q����=��Q?c��B�?xL��A����Hxg9n:�h4��6��޸��GvkwU����xd����-���i�ct�X������x�X�,§�@��,q��6�y!^�NST�,%<�} �d>�h1Q'��Ȉ$<B�ʝp�xȓ���Nl�@���?o��]��Қ����VC��Ռ��^��=)'�Q4�P#vd�"9C�)�-�1�,��qѤX���c��]�B����[8G�R~ KE���@�T3 �',�R���Ʈ5Q�K�L�ד@��)��Z���P�Ľ�5��p���8��!��r�X=F�K��>�ϋ�f` ��S8�0�����⌏C�c�'K^3A[Nr���^��  }�RL�F%�X+�vV`�[���v{c���Ӑ�4J+���c6@2+��<����K�7��չ�!�9��Cgg��쮱,A��aFO6�@Mft���e��"T1�������9/%Њ�>q�Xo�-\���>ݴa�$�B����J/~�5A��-��UxO�f�;�0�A@b�[�n1��^�,[�y�b����$��['��+���{�(I6o�+�)�yo��,�ڎZ�HPL[IP����rlśN����?_N�1�Q�`�(𝮔��n��/�j���v	��8���,7���7�_�����p���~��}�HZ�����>t5���ZoTUZ�UL�Et,�_%���@� ��D��&2�!���f��zB���Ʊ��t�WY�ĺZ����ϼ�~s ck*���-]�9e�Z��"|�[{�ߝ���=�#�K�&�dg7������DĻ�O���2��0�[����n�M��ѕ�d��~0�E�?�~S�k�ޥ�M�����@_�Ѵ)������qab(s�ls�tpDf��=yGZ�+-g8����u����؀�K����Ge#�l@`7���Ĝ��=�07P�񈬑�=`�~��P�Lyo������JRd�n5��n�r"։i�.�i`YɆ��X���!��K
��sp�|X�_�B����3�[�mg��[MU�ۥ�8�$a�7�K�0��I�n��"����>��2Q�h�6>X���Uvs]5��X�z�N����3��s�	�]�(�פ{{��/�	5��V�=��RHL�.?�Z��.�����2��痖Œ7[o�ZRZ�d0�/�
lA'�u�3���ʜ/NK�	��T��i������>���~�0�tGOj�e&����Er"u��b����R^����y:AKe£��A�٘��B�}�H2¾x�g5�����]�((5���٢�_|� �f��e���
��Eɲ� ��	bZ�i�qܩ���j��j��l�b?�2����,���n��J���������Ĝ�KW�f�`�T1��.̗Ý#��B_�\\�5+�;��� ��*������^�����&��@tJ�-M�xd{��]+&��gfGN[P	�-���+ݝ�3�o�kr��7q�R��MUֆ��Y>�vT]7���ԗk��T<�]�/V��
�z$��4�n,�c?\����R@�\�Ubk��&������Q��b�ݮ:�]��>A��{x���)�A�q�r��~�dߪ��`�@�u	��v��vm+����uL)ئf�2�l�-�/�D�<Z����3>y	<`�}��2��ٱ��+CJe��DLuI1�	rJ.�JK��柴5�8��8�<�}0�1<��'`"̺�l�[��t�)`;���1׫�&���u�b齅�=G���,��C�G�qX_j�u a����Cgiː](�����F���C���w^Ӑ���*�:C��8@�A�8��e㟵,�X����j���2%G>5p���|����̚��|S�>�D��v�n�Q��FԤ��觽ۙ�t�D��q��3�a�5f��� @%{5��2H�'�S���3$��q� �/�e�i�Қ���f��q�,diW��f�h�+ϻ���s&�Ƀ�$�UY0G~����d-6R��S�Žj�s߽� �>.����۪8r$�+�M����rc	|�sc[�>ҡ#sleZ1i,Xr���>�5���t�/�B��A�k|��i�������.X�8d����i��o�haE�[垮�@T�"!mh�Rm�y�NJ���Jb�K�b�ѳQ��PJ�\*y�gi|���\��n��Fݢ�K&���_Vר��[ZE<Jl�,�#K����Ȱ<�����n��I@ٔ����j�d���*V��r@_Kw���Ǥ?J`x�ߍ��QO���Pf1JV5���2jA��nݐ�Px���\@�������{�E�HJty(�ki��j�K�n}���` E#i����f�@����@`�|G�#�,��ɑ�����SwƑ����VlR�fR��R�&�4�O��сe�:9�[����k ��L�L�!�p�Ы��Ⱦ��T�u`b�<�ݭ�֡k/a��Vm'�宣�Ep��b!]����;�F�wS_����L�s�Q� "�|�W���0���a5!��c���O�[w_d8+�zj�mQ<o~�h�e~�2�rC����h�m��qm��7��\��QTi��;�v�&aLr1N~V�7`p�s�}=˶�k�lɶ��y86����5j��@6�;[]��<�ֆQ�]��jw�g夲��-�����nd�v]L��X�@E�a�;�ѻk^D�ld,��قC)U�v2�pg�N����YĞ�مγ���_s�@͗�I��Ĭ#�j��$� ����8Zy����``E�Y�n�I���2���1"^�޽��|�h�u�b�a7�Ԑ�����pIy�0����򟢠��j8�Lk�O�*w(���O�J)�$�:�a��ur���B�P�ۋ8��F�ǂ��ꇅi�87�Ɂ�AB��P:[>�a��9�3r��j�0�7 �4�e�&<��s΂�#��<�}[M!2:�P�!$-{~�|��Ʃ��:~����O�tKM<s:�?���85�*�+"����Y,��ӑf���Aw Ʒ`v�T=���3����p����bz);�}����#��Ea`��O��vz���h��M6��GoL�e&g�ikҵ��ow�:s�|�d��43E�^��h;�*��=�����gW��x��QF��<��|#M"����YL�5�������tvF/dJ����/Y�31������l��}�eL������&�+sL�|j��T%P�1�#śb�U,��Y��3C����;�U��ψj{ǟ�����ލ�[72��R�����M�e<G>�m27��b�ܾ%c���`�[���f+��1ZH�Wgh�xb�g�5+{����$���mmҁ��>���� �������W��%@�\�T�� Rٓ�.�	��BL��\G��e��N�q���#�(} �yΚ��C�w��fT/x��7�1K0%#B��%�Y�(��8�X�ˑ�
���71��k��� �Fev����(�3l��Z܀��A2��BMBВD��ʝ3MH]A�)53��8rj�͐pn���?�I������:�G���V Y�)rGg��>���o/���d��9��RO�@Ų�a������d�2p7w�Ϲ��?d�	��jF�E���%�7�w��I��
��Ŏ��Ӳc��1b7�{���ؽ�;?��v$�h�
P�#��y$��=`�s*8O�ж$IF�pc؜`���3��"�a�~|�=P���LL4@�� �8-[O�%���G�+K�Pvp$EF��/<`��9�]bVL��G�k�/ �~o���Wλ.:X����=4�ȁ�Lpq���BǺ�k��$�h��1H=�X3`��){q)Jꜷ�}0Ks"zؚh���|;	�[�z~�'�P}��N=AH�I�\��y��8"r�)1a ?DQ�a!VX/ɒ�#���G�����9��ϻ���S|�[��0-�ܲ�A#F�o��,ܶ6T�4�	���m�z�`�l�,�) ��׵D�e��-�xZ@�:�����`m5�=zoT;����c�����.9���n[�dy��H���_�&��QN�3��0�%1bŰ��Vb+D��9�=}7�oP��^NA�mBnolOyk��l�	�T>q.���Y(���b�wqQ�ګ�s��fl�C؋q'A�K4{H'���������Ԅ��N����~��Ч>�c_P������^^�Eb:��IB�\�,3GZ��X�C���W�)GM����XT��QE�+���U��5�aw�6	�WS�	�����s�/f<�ݻ�KX�>]w�(
TȖ��x��e�i�շ:�u��w��1�f�KSD�%CE�q+$��n��$3�����i��6K���{�ꛍ:��3��c"��� �`�S�"���qC¦�O��3]u\��`eyԤ;��s��!(��o����B����&9NI@�ܭYc�.NE�V�O��%!d�t-.k��!o^'�����,�FANNȦ�J�
T`<�OIkԓ�#?>�)���p+\^�_��Q���� �v����؏�N�����%A�VK�X��*/��3jG�FH�E�,cc($���/��T��E5q2�<�u�o�K
��);�R���0��@=�P������S�Q��ޚMC�O��ʆ��E Ë�̬^��f�(�+nAp�=�{Wm����U��W���f+*0��B��멗�%��G���)s[�R��$��l��7�0I���/,ZbBg����B�D_�8:5��d�~�:����A�i<�9Qb:��V��|s�i�B]�s�W��~@p�#]��@�9.��E	�'�n8q	�^�a1GY�`�ܧ���@gܹ4g���f��2^,:^SZ��3�H�;�0���UP����=fO�M�F�ʐ��7�P��i�S���=�Y��+�WϚ��,��͑���h���JԶ�m9l�u�>H�Q����3`M�p2���	+��#a,�8#���6�{�1ٝ4$/U[�Ǔc%"ƾ�UTk��C6�9�I�сڙ�zuf�U(q��Z�&����JI}�U�ÇR�B�������N���nۋ�5m'd���B��\��sXU%��:l����L�R��M�a�x���p*�'QS��z�ᶆ���}��j�>Jd��њ�!s��$�p>��%S��׊ߛ��o���#�x�J���p�"��%?q������'��� 5X��mW��c֚��/J5p �x��[�q"�h�^����OE���O�qb���O�7������}�@�=�cM:Y�4���+�'��@Eu�߲x��k�bvѶ�&��U�s�I�s��jΗ�_�6�qư�W�!?>����l�՜�ƈ�W'D��x�t,��<���ƺ��fH��=�k]��V�F �A� �Y�8
h�u�"�H���F�R�xq_!�F�I�������M�ܣ�'8��=]]���u����ձg8�b`&�b��^�y�h[�����	49Ay+ֻ�Oc/$5�˺-�5�7#�}Lt�M��["2A@�l��!���X����r?�k�ȯ�a@��3�?��h�c�y��f���z�}�4a������DGC�ViF��J���w�䀕H�:�D�a��IV�	a;;�)����i|��PFxr�B3�Le�z[Vh�|n�%�T�8�L
�;�5��BF�J��M��n�lT��m��������pҤH�qr4�D��Ņt�@��}Y[�	wO���F��&E���?g��?�eV���!�g��W�|G���}�'l�������s,M�jyh8V���<r�4jE3:f(V׆'�鹱G!���ON6%Zi��D���]f+:|�c]��3���A1��{Mzs7�׼\;1!�!%'KD/�����ؓhBk�v�ʚyt7��W��#�C��g��������"�u�v�xh��U.f��m����<#z���R`���;���f�A#F�[�`�C�*�~�J����13ƫ~i*�FO�Չ�z�͜:������]�22�w�_�D�����Q�F�m��]��ǥ�/��_d���o& ������y�4�V)w]i�{�G��'�ˠK��W_.G��d��H�\�6���w�|]dʼԗ���ަ��Ȗ������\7�rI��8�-�]��<�@I7���(r��2�����Q�[�\�%���Z��5�0���*�&KC�O�W�mLZ.m��.e	u���WE<D����мǊ���������RCb9�D7jD�D*\`�DS�<�?~f�O��;eQ6X��``�Ʈs{�����<BM�����]ۈ�<��^�<t-P_��҉�%�6A�hE�Ʀ0H��Q��|�QXѢ���|ao�Y?X�ӝ��>;e�H݇N�'����0����׷�l���.�r��z���VO�G�P��`��ݤt��%�]j�ٽ��[(\'�H�_l�
���jR�5�La7��	��S�.��x6z��c�dt���A㟸O�O/�;�5rr�ﾎ�g5��9�!ų�f���B�3zr��ɭ.��9�rh9ͮ�`3����E�\�$�$���3)9�^�۟���ݽ�@��r�
���-���x�^7d馶@��+���s\u�E����Z!��Lm,ҍ-V̓Lf�uѤ./�g���N�	��
D�_@/Ϊ�=�ۤ+�@N7UL�*H�W���A���LoЊy�<1`�g;���j'&Qmqug�YO��9L�A�@]�)uv�~~�d��+q�Ԋ�h�~�<v?��4�Z�z�%��г�c=��'�5�<�b'���`)���H�a���^N��x���2�� {��������tY����i��-�e=�Z�g�x��h�i��3���W%=���}�'ݮ(���/?PV����Lz:f���y|�ő�̀�.-����@�Y>���6���R�@e��⯼$�w�L)�~�FEܝj����6�=$����Y�2Ld��_�Ü��~nd&�'FN*�~����>���6	e�E�=wn���Ys~���3һ|�4�E}�5V1̷�"�����A�R�r�eH���ff���4F?����w�-I��_��@�_
�p�t��M�W_�J��Z�L�ڍ"*�Ɉ��\���K$|~��b���[�
ՙ�孟��T�Q_�7��:�J�ү�R�ŧ���^�m��FP�����.��w�C8���4��M�d�7��?�ּ9k�H�jKU�{��H��E���R�\F�\ ��z�b�UJ(�UHw{֍�1B]�=�Q��TH�>�'h� ��
aY�_I�㫈�W,�ڢ�rN�Mx�Ԓ�����!zt'� b�mI�D��R�Q������/�}�����HC�0c�6�ԢT�R�/:����1"J��!D���~-f-���2a�f]���]�W���p #�x��#'GJ �ŶD�r���Μn(�r=-��|���i���P�8��9�Lm�{���gN�U8@� 4PE<�� `��y� �áL��jS&�w��Oʚ@4\MqZ~7�	��Z�(���hd���<v��|����P��a��4Ώ�H�0s�ja��`Gj-�����П{��TF#�ʔ�4�CEH΍�/���tʌ���߁�7�P�1�W���I*�~���'�c�j��8����L
JE��λ(^	��@����O�(p7�V�x�z�f;�RQ��EJ[�'��	��L4��%���bNB�&b}.ܼO����2wu��a�5�a썎�茋�x�Y��l� D�~�~L�gydcx�؈W�"��AyN4�%®ֿ����a7LO��l�-k��ݔ<��[�18�駌�j��k���(|��=�Pw�v���\��͛�F��1-Na�z�8`̴���W9�O���0�W}�
�[T����wyT���^�G-���ѣ��c���.��"ךU��N��� M}��mC@M��[��� ���{��c�}�H��/^!+��D�U�2��!��1����x`�h�[��Y��v|$'�-3w��j�L���~���������,b¢=ΎW"t�/3����+��=�+�Rr�6fD�tv��Z����U�,�� �h�����٧�1m����Ow�I�tEh?�wRw�k�RrIѰ�����Be��[Y/������{5��[���nF���eWs�<M<���$ɻ�V��p��`�mF���0���k{k���B9F��I3Y�����;sE;�I�5n,(�ΆC�/�(v}{���Z�t�#���d8?�����l[��,V���TH��6�7L�in�6���Mv����@�b�P�`�?��#�e&Y�RR�z�[�1��+���e*�OuM�e�,�ֹ0~�%�V�?�^�C�<�PY�rܑhW$�n�x~���I����pB>���db񳺱�]��i�ꢒ�Ѣ�"s�F���)�Խ�h�)���ek��Cߌ_C�28���@��Ӯ+vߏD���^���"2*�ա�7��g�Q���4k!M��u>�Aŀb2'�qw���:�K�Ti�EÞzå�����C���T˰��6�}��󬹌l�{��T�^�3��HRq⮠#���������H2��`�K%U��+�Cg}�n!	p�3�y ����&T���+Ɉ�b����W�\,�V�ef%��뗆ݰս��ݣi<��������\��a�9��)mo��bN ¹�;H�'�� ��|��"��l�4
�����x�A�g2���kC;h�w�=��0���� �K����q)��p�sC��@Ϙ���e���g� �,���U�bO"M
_�<���^=�Ѽ��7j�t"�5�<�5��ܪ��]�X3G��*d��M@Qç8�ߣ�k�Yߡt]�i��zg{~��x��j���df��F���W3�r�vǕO�������+�z�:�E�I^gŀ�L�Y���Ċ��G�`��Yy�iQ���S�lP��_QY�_u��-/
O�?w޲�
`�k��Υ-m؊�=ii՜a��x�?���ZC@e�T����1!r�S�5	u���dҐP���:�o(����ܭ��^ _�Zk��M+��"��#��^��t?��+�h������q�E�:�%3^���q����7���(��|o����N�S(�*�&8�F�DF=b~:@�۲3-�^��)�\�I���I�T��x3dF18q�<�V��e���Q��]�N�"��S1I)� yx;L=
��v%����l��]-�j�^v��L���^��]r"KGG
��-T�TR �Wg��_R�?���()������2s�d8�3�I`���E�f`�aQ�
���G%�Kw$�x@5��.7�@Px�I�3sx��K��Lzn�QS�"&�L���#Ip��?1}j�>�h�U���:ҭ4� i���ܮ38����������=�4���6�Ѝ�	gШL�n���\X�f����𚧘jl�9 Tn�t�A�V;ˎ�9cg��K�����w��\����n�O:�&y�&=+��27���M�k�bF+n<���%9G�pE���p���,�p����u����*Mr躚�բ撁i"u~ |���F���4�؟P)�<�&J���0&��8J
:����3����������6��������4!�')Ѓ�̃���h����K�.h���	�l3-H���w�ǉ̚�]�h/�/0彎b��t�VP�A�kx�ªT=���f�ɪ���Wd�s׳���*L63�. M+Ȗ>�m����1$��.�F�Ń��p��۬�@�[����qp/�9�����ƞ�8�r_8V\o����Α�ް����L��go)�#dO����Wz�y.1�MX�����z�����&c�#�k@0Ty��>g�q�������@��4m�q�p��y�7<�;CL��-%A��&�Qda@4oXB7H��8G��wd�[p�#l�ܪ�6�nb�����8UbSX�|;��R�A;B�b��˩������(y�t�����^˵<SDowjt�zM6�\�<j?�̎��
�7��y�%}��^��؜��냻l=��1�'���Z��5paŖ\�CG=�vdіY��������?5����I�����'�})H�PG�.M��).�J?ݟ�_z;�ߓn��Z
�D�(=�wM.a�m>.w��{�4l��8[ �?�}ŷU�Q3fFW/�ؼ6~�F�Jt�(��8���Z�ɓV�Ú�ŕ��o�T�]�і/+z,*<������2���ZdXρ�d?����[OF������ǿ�J�wrKxR3Oa��U�i,;���5��� ���#�Y��m�w0c{XN����E"����ѲYg�c��������еk�ѷ]�C��%�+�\�${J푚&�f���_�J�1�(����Փ'�Ƈ��)�uS�6�g���,�� ���ŒL��mX�����;jR9Fm��_������A��-ۻ)��B�8�xh�@8��c-k��Kv%И_�6�pU���vT�c;v6\.ޅ��ePھK
}���x�DBg���خ+A����*�L���X����Sr\�nqE��Q�b�aYrys���7�Py�RDZ�1���t;F�Q��D0��n�xJ@�JmN%��(0ֽ P0�}�f�N�.�d�Dδޝ;,�P��!��rm�ȘXgO
���ψ�A��?̨�����ƉjO��Y���S�����MyT��X�Źi��0�����X��O#�|Yre���GH��}���X�V9m:��]#��V��?��tx�$�����#,1qhSc����,�q$�Q��]rsRp���Һ����ࢉ�Z��%��Q�]]������$k /md_s��6"�|]̜l���&���+F�����j2u�nU�!O��b^va=���S68Z^���w@cr��vo�����#t�4���V1y
�NJY����A֎$�\4*����T���}I8�0�&�{�0�.D���W%՜��~�ܯ	jm3O:��A��f�����V����`��z=��B<q�<�`mD�(�?��y)�}�|39��"����B�X���w��!I�����?ȸ��pm��^-��g��_*��r�LD���׎�6+^��ٹ�S���1�j�۬H;9Y�'=�y���kL���嬉��P�nD��ߐI,���	Z���Lp��0���"l|�ŝ����?G��]��xyS.��?�gi͕��2��.�R(u�/�>I��Y&��NA7�Q	ؤ�l]�e����.S��W�3n�tt����5���.�
g�N���M��}����кU �.a�P^�5�[��Ϧv�0&`�����}=4Wdio�K��vd�M$�h�j�FV.���B>����|k��ч�|���*��n��`ޘ<`;�i&P�Y��^�Xjz��V&��p�(y�;�k.x��I1�#�Ma,aF��A��RF`>͇�R]�u����A]�P���E��|&d�����]�JY�U�@ueCuA�b��@ld��8t��mƏލΛ����Ҹ\�����Ő�N�*p��N��L�`��xw.��� �����w8������w�]��d�E��l&1���,e��]�z�g��0ۡ�|.�� ҩ$�N�j~<�������������]L�gX��w$ñ����~��C�|D�����M^��� VA�������vh�;�=P��#f��||��]��+Jnf�0���Q����(Q0u'��œ	�ǅ��en������{T�;�ы���菾��ʲ~��|���&7՟�گ�ɶ��f��{|�e3�D�^�F�Q�n�fN�8�b��'X%�jD@SmѾ"�򏐟1%x���W�&��=������q�@�����F^C{���	����D���a�G�f^�*�:�X4���3��q	@3������gQ�tn����B��P�����.Rt���t+o」Q���RB҆�~�ZG���iR5�����5�UhCI�I�frxz����ח����Z�4�=�&�8{�$1q�b�M���xjM3�W!�lFfN��o��D�z�nV�	q�����00n�"1(��R�<�������v8o��
xր̀�9P��b�&<���6ڽ�f{|%�5�1�ٕ��P�[}	�m��u�W`H�,�	x7�Q����h*��/䬣����˯�����2Û�N�'AN���*0�k�&X�_���81B.�T/����x�7��w3"M.�6�V؞�.��d�&y?���f��pR��8���@߸�)��>���IY�-/#~'� c�˼4Bk�"y�l���	�%	�CdcS���#T��ũ�gr%N�S&i-����>�V:�*0�k�R9Z����'qq�bu�sM�R�`�F�K4��<]p�3�RLƱ?��*��m�m��h������'_-N;�7+U p��$���X�"(W"�rn-�/5�?���Tt<4� �&��'�I]xP0�y�~7�S#v!�\�2њ�����VK��f���tr+>l姬CK"	n�~I�걃�Dw��IVzӅr��{!��) ����㌤n8�u6!�/����C�����QSa��FΓ�w��^$�Kw�[00>�������N��{.+R.��	�m�0��4���8�!����9d����(�Z�W�q4F��s�e��aTWW@H<����"ܨ�c�W�~�@�`�;�����,�����!��+Ғg��ڶ�q�H�D��������cԑ}\lp�qڄ28��N9�/�'�[�S��ܐ?⧾���y��@�&Mt���KN]LC��jw(�C��|7w��\�	&13,���@'M�t��Q#�FR�\Ժ)�����bt�"��.�ǈ��h b��a/����L_c�v�M�oi�0�gnD��37=ĄG8�c��6���M�!���0�F+�J��3�-�ҨG�AIt����i-d�W���m�"m�O��v���&�ͷ�(nY�9��@>X�M��)���騏��0�J�H�(<EJ���>L��=��G.��N�Q��>�ﺁR޷Y $����Z��9Ҧ@��A�Y�*��H���n��$I�Y���XQ�8�ڐ��Řn���B�Z�W�J6�?}���!|���I��7Dw�g���*�O���Bd�沎��Q6ރ��Y󭕜��BX�4�,�_��¾U�/�Q\��I-�M����ZF i�\���I��ۃG~_�>J,R�,��li���5�:9sVs����L��p(Rg���U։�r��%s�sT�2���%wu���Z^��9%ڶ�h��k�<�8��--5���e�N�H6yi�R�#l����fe��|�>ȥ��]�F¡@��<z$���Ҡú���zpA*�}�Ȑ�?�$��8Ч�����1�1�~��:e �, �����IA�ޠ�bXW���i��������Ij{��6��}��ė�ׁ�Vlz��I���/|ih ���0=�"�/�CfU�}&�������D�$��$�컡�S`c���Щ�s��<?~r�|���ꚝ�N�ޓ��������۽j5���g���檐��	m%dB	4��-��'i�@���;������TԜ�����_��z�M/:�Z�����"��}�����U5;��+�����	��iTkN�ۆE���sG�V��*�T�N��t�<���l��r2( �r;�nM ��^'�ˬ?���l�Flj��=�o��E �A�k׷+�1l��LOC;���k8�P��P<W`����T[�tN�\o1�|���@��gѝTc�$1�p� 4��kt����^��ƹ*+�e`:I�H��$-��dF���r�����m��'�J�:�0�з������&�5�I�ւ��t�?�V�J;�03����JM���Lh'��E"�y�O��8#O~$g��r��-¯��s�(�����Ɵ0��{qr�O�!];5>l��Mk7�A"�S�E%[L�ڋ%&�~ ��p��%8�Z��L�MZQ"�nFk����F2�voӵ5_:{��0A���S���~X�u��x#%:�^=�3���G��b��/��(�r�EE���)g�U�K��F�Y���X?�ꟁ�}o�O�[$�*SlFV�I~�XfS�:���⟾9N��h�C���1�޾���[=������ �+�1ø�ˊ���ލX8��V��(?]��yǝ��U�_\��֫��;8n#�[�ϛ0�#A+�\���9����z#��|��N5֣Qᆋ���cY֛t¿)×H���� },�2��u/s�Yc3�w�������>��S��J��w)w?���dT���F~�t�v(aO�\7Q�wP��O�!�GWfV'��n����qƼ�7�j�3aÐ�8wYY�����Pz�;�ʣ:��օ� �'i`J��]�V1ޠӗF9lE��P�b�1l���?S�~O��Lq���T�&�U��ĕ����1�=o�6ѷP���T��R~�aq��!��{�
©��F2�[��Y�i<t�%��n6�;A#e7w��_ 2�s�=י������-�}5�٦F|���=�����P��K�%�_�^*�K��҄�	�-���L�<`���r2ӈ`y[�N�tVЄ�I��w���?���N�a���-(I��� ���z������.�~�
ds�o%�(k�g�� ��r�*�d���_�)��`j�2YI6V���كL�	"�J�/�:�=�70fc�	"�i���t��i+�G��#���v!��I���-��e�����u�a><DU&��8��_�t����E�aPJo����w��"��l3�+a��!�X; 6��Jy�87�#�̝� ���*�#䬋D8�2JAn;hQ�����M�fSI���.��>�&2�#4�K��O��:��pm~�~A�tj�U$��Ǫ[Q嗳ǫ/�T����E̱?E�!�I�!�����0�=�ks�ɋ��1}ͬ�l���v��i�Ϛ<RRF6�~��4ۑdn�� PL ��������<� &�7�X^Y�;�e�9[?�#ݗ1��ڳCIJj����=�ե�uP|��s�R�fDn
�;���8�j�#tt��j&:�w�0��FP�WKVr�,�����\�=��i����ɘ��t�������M]��.z�K��s�%�٩#���Q'�x�:O]�c�ID��s��cG�F��y�6N�?n��K��/`!���^�dC�2q��sk�[�(C��ɺ����klF�	"��IK����3��؍�'����w�������8a	���jsb��5ٹ���&��\~���-�j����E�7�EHm�����}�d�i �*g@�(��#�(���#C��>���p�9!n��H,}�V{V}h�i.�Q><$甋�o�c�L�H�M�Z���B��R@�)��C���2��	�_�1DS�&���I.��J)���7�4߷�d�������izMm�����	�]ҍ��그��`��{`��Ze�;,Ը}�W� }C�؅�	E!�kG��ZcD+��dltLyY朗�e��GJ��/�x�2?S��MX_�L2��O�/)���I.��ȵd7�r���X �ռ�G������]�<w���k�Ra�Q?SMN��#e�}I�m��v���I��F�A�go��N�GC?��� =:�C1?� .�U�(7�b�#uFZ�wu���ބ�F�'�������C�e��S؈�e��o=?|S�I�\����g3V���� y��Z10ݽ��P�/�Hj�Z�E���О:��W
)y�0�yT�K3��0�tO�� �a�� k�t��ԫ���*��k{��5�ޫ
��`�+�F߻������f�|�!=�%򱝬a�+um�:��J��ȃ�Kڌ�R��;k�u���9L�S�@�yh!��sQ� >���@_45� ˯.hRAk�V\K��$�j�ӯ�\ %�0��Vr�U�_zkV��"͋B_>��+��!�pڸswóK[sg�;�:YR fF$K�Rqm�5]��$l�ی����ax��>s�?�o}�#m �~��4�nak��N?��C�y�Z�_NAU�#��jG�	
��J��ϝ�9��#̦����#!��N��*���,�ّ�����]6�K��}�j���.��n��m
J�}8^p#;��*R����HJ�aY�G� �p��ӂǣA"�5�W���t*S`�K��C2/x�p��Ԇ���*�%D1�y�JjA?����I05�^S��5_�Y�]���q�+���`�\E|�-ɚ1�\
&�\F���`6��l����'	w��F�}�-G8QejV�vd�U!o���x��i/�W��W�,a;�����0�ޥ�v�NI;l�ˈ�~���Ӏ,���4����2�$Ȕn{�?!,�� ���Q�Tm�R���H?
ՠ� d��?2#��l���'T���;�~]�Rg��\U-֬�������9w���2O�����X�uVb�Xו�끳P�Z��� �/�e< �6mE(��am/��)Ŀ/ї�nN��������5�,��Q]}�p���o��fѮ֑��Zj�|��ᮝ��0�_�O7����'����s:P]���bE�'b]�1�b|aY����lj�tM�^)��F7�](LƆ-�'�
�솟"��g5ᇥ	A��=�?��ط�K�iXT���A���+/��L𳜣;ͺ�a)Ⱥ���A#c���B�g[�{���W�
s|�f:&~�=���	�����}���d��ݞ���-b�N�ʆ�L���8s�
q�������2���T�P�V"�)NBP��E�]և:��zT��t����M����l�1вV�TB�4D���{���ů�g�9�@	��nvzJ�n��C@�9��2�� 6U��c�����)k��18P�5��=*��iF���t,+|�"4�Y���h�����;J��1ͣ�Q�*�`��b��3�j�ω�	0�5�S��t�����8��uǘ����NNB;���7�C5�y@��K������ A��D#�$܋Jݸ�Ɇ@Ӣ$�C���?�86>[�ZVP�;�*̠F�GW|�4�e��I�&,&=���0<䫧��$��ѵ�U�3���i>�6�9[?�8[)��a|�t,c�R�@�Ͱ�c�{D2��XK͊)�~��#��k���1}�J~�6�H\�U�v��*�mk�-�����1��PWw�\�:[ס�Fyb���[u�G':�\M6C�!�b��[Vz�#����G&Di�X�$*<V�CABMѫ�Z1R}'��yݚ?ҽ����F�hzQ\��tuz쫥/��G�:N��T�ۥGY��[�V��5kT ���CR��qA���:��o�/C׶��Id�m*FA��P5���q�G����daAد�B������Z	:{<��C3*��R��-~�B��!a�or����{|5�o/7�X��t�֑o�N� �*����4��Y���;����4��Ɣz
N1�9�:e�Sv� �:����%��>rY�����Xc�?W�U�6s �gB��(u>�P�
�P��2�`�␶pqsmt�^"��m����s*��������V�*֠��n���g3������j�F�� �;u�F��|��eNH=��� ���� �6&j4q�(����L>u�p˓��%�vߨ�s��T���2D����������,���]F�����8� ���_�7kj'l
N���A�B�[0� ½�B��d�v���5"{�Nm��V�'�?�1$��hF(���la�]�3����t	&,D�&\T�����r�VF�ea(6]?�ˤ���]���%W�8�X�I��"��'m����D@�J ���;nTF�C�pV�/,o��w9_��s�k�ۂv���`��e-���Ao~F{u�{q��|P�I�Z�ey.���=�I�-�n�>������.J�E%�j�I/�/m����OH�8�t�F����*^nLe*`��i��,��o�;h��2�ߣa��m��Q}��6M�󏣡�G6�=� #�B�'�Y�D���P5�+�����)�,ͤQ��:b��Y���O��AWh������^M�Ar��G��|Ё���E���Ɣ�X��lS/�$D�¿���2Z����4(�yE5��F8���Q_�&	v70Y��&���<d�i/6��ic�5�,;,��/�����};�dd��O�1d����h�r�{���r��]�S�vIOZ��/�k�=i��50To�~m"�*��(A	�U��яI�j3�-m|�p��w���1������UK���X{�4q�"Hp��q2���O��7����x��z^�+�ᵄ3��Z�l&-[�_0���Nz���^�8��qm���O�7>�P�(�y��:4��͎rnS۠�`tȚ�{�ŕ��HkhB4��SC!��2ev���^�R�o����}��j��;�Z	Iw��яW�b�Zc�.�;jTW&�l�R?���f�s;��V4)r�����O���+�f��&5"j�ԥL?M��(!����P�rW��~����)����9��a�B��3�3�`�tM��?:sUK�ה�_��L#ܝB�J���҄<��R3�.���V��z�_��-�z�U�����lʎ��9�$���^I�i�?���j��,V�}���}*|D���P��.�.#��x�a,���d�4�j\S*Ƚ.K( 0�mO-���Nl���N8~��1dq�ҍK�[m_�������)���.u�=-�4���Q\��������������i�m����ؽ0�}E���5X�	~M���G��y �z��W�H�4�
�%�?���ׇ]��|8X���i�쇔 MU�C_= T�C]������InB&L�O�"���X4�zX����ѩi�}m0~2g=�7���rF����ヲp�;���Y����(����_��__��"5k��}��B��������A�"������e��8�IT�d�N�P���ä/�	O�+~�Mu۩	�֢@�I#M��P<$�:q�/m4��]������4�����6D�Ѣ�1.���9jH2+'�/�8���j�Dm�#�%��g�����^�X'��ᱵ��pF'�+g&�/� 6-�8J	(�1(~�7v̳1T ���
��lC��?�y.�ҒJf���5v�8�rkfS��bͣ���z��d{��;��3^4^�����F�0�|`�	�mB���^��Sk�/a��$G����<�H�|��|��
��~��Q�1����ړ ���4ꇻ$U���y�����&)c��(�o�V*ν F�,�&�������q� ��z���ّj��N�q��������xtcgԫ:�$��3����b��u����I.q���m9�y+w����Y��7�����	���㩞izI�r1y��M�� �o�.ΐ��-r��@M9�K@Ny��;W�pc��'�B^�o��&���g�Ʀ�j��07P�leSvǧ���X���K�WY,M���d�"���\�`��>�(H&�u, ���<��,��&��'vI��o�Ib�#�����!Tg����KYi�p�,��Z@M�H����*��CńB��OH�[tjF�v��Y���r�^�B_�LH�L}��H�	���ؠ�)
W${[�A6�%� ��j��)�Li�u�۝�;�S$���Ekk��RK�.$�� ������!��ҹ=M{��5�_<�ܗ�/��YT���bܘEE��tX��a���g�~pf]}>´��Wu�;I�\�Ͱv�!x�^z�!UЩ��� &���%ȍ�����xe��XR�0��_�72H����dM�gҊo���7��%���b�3��
G��!�V�4.�T���jP�-5{~oܼ�BdIg���$Pk0k�O��y}^8��hڗ�S�� ��N*7������l�x��:9�˘��{������| �2L�������&@�#ms�i�Cƨ@�������ʍ�q;/���Wg�+�vu���Y��"�ji|�g�D��j��(��$Jd�m���؁!���7[|C	���K0��N��h#Hص�uh��_�F�@-mhŘ�A�o���y݂(�i�cx�~ϴG��7��[X�s��H�md�p1.D}ۭ@��x$'�F�\02uG>�Fd}k+�s�z=/R�֬{sI�"�	Va5R����1-(-T�Ѭ�5_�����!8�#3��ON�s9Զ&Ԩ䰒(�hJ `�OX!5�=B�
L{�gzՋMYMdp� ��x4��ۖ�h�2�	�R�xy�|!H���wl��b�ʕ�l���ސG !is)��j/��7Q#�!u-�}����.&E�WH!�R��%'��d�`��� ��nv����� �ݡ�Sk���a!M>I�:vfV�9��@��������i����*��.V{:��{��*k糞�0��8��1\�f��Q�4�;�޻�V�����=��kef!�뤻@���cP�αh����O-���Tj�'�Z ȋ��q��6�&\PR4;e��t��X�����E�n�j���KT>��� �,qT���q_U��}�`/��	��>��'?I��ٓ��.g�[!^D̖e��>$�ڲ�KF<|�e �3�b�:)�Ԯ��� ���i����V����J�G:�����f<�B��?�k�;~<��I��3��_5h&X��~��9{L������b+�[;݁ě��$TR	��$Yʝ�:�F]�!�
ϓ���:�k���lջ�#Į����+K��*�)c0�pj�e6�=o�#����H$bfO��6x�p����m)GV�σ��߻���$�N�^��
VT�����e��)�X�D���"�6��<�O¤,?�� ���,�~Il5W� O�?b�)&ú]8
��B�y��m�$���JL�1̊40������^&z3��N���k'�c�뀔@D:Xb*j0O���R |^��IcK�*��z6��rL�w�F1ђ�
�"����n���框���\΃�������#tu���M5A�I� �n��f|��O�[��t���
~;W=`P����^T�R���$���
��r �#��������a�k�@�?��F��s�+�!`�6aڹ�f44�G���U�y�d���I�Q��`Ј�-*�v�I5#�E%����=-fo�!�g5!ˠ ��7�5?�}.���+�zXg(Q�AF(�k�س�D�F�0}��{C��J�ώS(����ҩ�]Ixy�ǭ�J��p%o]�#�gu{0Lw�fG7j��]�z�a�i=�K��W���K�4Mp���pR�P��ovPN�9+�έ�@_?���F�k�B���ZTWE���� ����kQ���TԻ1��)>÷���/d�0�ۀ,�u���.���0��Nm��s8��,�TK���裡%ª+��;d݆W�G��a��� �e��j���+�O60�hG/�@p�9g�]���!�s���o���n��zϜ�ȅ;9�h�q�T�c6�h�ǀe��I����5c�Z��dl�s�Uh�O�7"�����N�d����$S�׭#�|8��u� ���/����'C}r���jJ3їL�·,�$4}:t8N�țH����a��B8��Ji�!�Я�YxQfI�g@�浵�H�`�#�����ڄ���8�&�9l�Ь�������u�9P?�%#��/��&�|O9ժy�ވ���x���m ǘ"�Y�O��+�������y�B&�����z�%�X���a����OA8�̸�8(��UB�{����0O���1R(�a���rUta�*7�!)��.�ִ��C��G�ܓK�FV����]E
�ŏV���;��3>���ZY�*#��-AO��R�|��б,,3J���b�h�\�p�]q���sů*	��!�-P�z���)�#HwO�z����K��<�s�8�ڞI�n4GZM
+�+�`�_�0��$�#5C���ۮ����m̚W�M�A��WYWE]��ق�hx�̒T|6����HGgrS�t���^�H�p'6P�R�~}�F2ݵ0H�w��ƔIj�e�2|6�J%ed`L�\�r��Y���چ���͇(g7KOq[1J�8Bn��X]�M����V���&xٮ��/��\��;������%�yJ6�^C)�㹈��8!]l�1Eꢷ�:��X��,AoB�yHۜ`���uh���(Rء�S	�ы�^�\�x�v��������!	4][0�9��s��CO�O!���/d%���
���*���j��s~M��b��x��[m�9��0�!��w̱N��`��4�2�|��'����*�gq�aqԝ�T:��2�5��89��D�$,����F��AW�&$�u]�^&�uv���1���k�j���������z[�T�����,d7G� Ke}��%�/�F���e�/+���{ ,�����u��_|���a��X�\�!4�!�L?�d8i���![y@�4����;�C�LC"/�y�H5_�1	�)��$������'*$�|޶c8hF|x/<B�]�g�4~h7�4���.!�5����w2]z��F0D��٩M�����\8����c�uZ�W
�M�^����t�>8�?YT6!���b&��+<m�0�0��Ϙ?�6�?]��R�lŋ�"�B"�T�J=,�E��'�Ǚ/�`/��҈�:�+aŘ��MIz��j2��;��C��e5���vF�㧄�.���J8^ *����:�^G��3'�k4���5^�f~L�J��Y��cՉ0"��e�f�X3藘�3���Xч��!��-��_�K��������:�0-'�C�?������3-n�/�F���:�-3i\0�9̖r��M�CAm�F�nj��L�y���*խ[�Oo��<��Ka!�y���Q�bY��Y�AT^4���6����Fm�H�3�^"t�q���'H�w 5���7Y�0�F�:�� �Yټ_{�4?���������������Z�*|CR�Ӟυ�[m�+as�)��E	xե��=��;݄�%�Z�EA����O��W�kE� V�д�'/��x ��(�ә��,=�|PM��#c.)%"PUMX=Kxf�R�!_�m��U��!I�dX
�	~�����+�\�V]�cJ,�bn���U�*�隆�y?�F�9������v&������-�=k��*\�_I��b�ĭc ⥲��4j��W�-`#��uܹϋ�,��:�?� a���,�?k�]��Ako���gF�� ~zMv�ʳP�P���-0���X�PG휬�_N$堘~O��r3�hze�E.�M�c+E����є���<~�$k��c̓���� �S"���k6Wî�1ˎ�HT��[�d.��$B%���N�is:Hg:��z| �j�(SB��{��4K����@�S/��2����wk3�?��u?v����ɀ_�����JY��-��}^H2Л�뱢�u��fE���)��S�-r�����獕��X�퀎u;�0"if)�gǺ�d#��CjD���1%x1�yZ��-���/�I4{O�Ҥ��_���?@㹬#>T�ݿ��J�j("S�rW�c�Q�|����e�CX��0
��%%�ޖ	�y�"�8 ]���~4�UeAy�XW��/��S�w7�'1f�P1�yoQ���j���+2�j�Ց�`����j��ۄ�q��)(�����ι�O����7�[	�f2�Sd<*�a����l�� ����%IغE�#�
�赊�xGG�%Gu���������a{5gDZ��!��Tx�;�nE����1tl|�I@���n ݍ�Aεޓ%dj{q���3���u���s�4s\!	��o����b�Un�8H'\B�V�� 6L��s��d�
�X��.����F�Bh��"WW٨jӭ8����Ģ�]f<W���3�;�$�O5����9k[ɲ����/�P��HHP��t�9� �Jl���Vבb�m�[iն��
j:���b������$(���-7���8�t�>6y{������� ]0G��"d(�|�@|�S��T�a5�d,��܀Җy	-쭠|u�s�=��w�mk�Mͱ��׵���_��ٳi<�6� l�%��	���'��h�
`��[�o͗-�2�>�����:b���n��T̔R��q[	�s
K���R���R��b�O!�I��@uy;�Tv���Z��(�E�6n%�Y�i�����*�tކ���ĕYK+������Uv
���xe��b<[w�?,���/��l`�<�7�; � ���8��a��h���j�^�����z��)�:���4b���-��z��������n�p/�Q�#����������9�>�s?�Qt�ˡ��W��B���L?;v>���uɴ�G����Y�퉨��u	E��,q�˖.K���m7��sҮz~)@0�dt3@&)�Qό��պC�Y�J�e�R]գIaBK3��������Q+o����~Dl�j�N
ظb��kbak��nU5�Z���h��W:�Ɏ�����`�Ol{�P���M?F�$���`����C�S��}S���`* �0��76�k��%��5�U�p=a;*V��N*��l]@��7z���o��5��@�����A�JQ��(. � �'���v��Ex��84�Ӎ���>�.2�p�.zĐ�����)��سdt�xHG�`�Ue"&��CWC�(��EL�BS$�B�;��D�A�zJ{@]c=��{N��Y�M����l�^�?ɟ�P�&�	.N"���9�N�,�QMZ�u5D�m�z�[�,�F������X�ʕ4��K�ޠ_A<����W%���e)��X���O��e0�Di9q%P\I~_�N��U�X}^HuRT�ᛱ"���-��pi(J�>����i�uT���!�YzIO �U~
��������� B�̿z��j[Վ&��s��?}�M��A/`�9�p��eCX}���q6�l���(���sH�:���u��#?A�eX��M����)�H��4AJy˕�� �;�uZi�@�f�ߢ�p�2Υ�s�0�YE5~=�+ES��:�2�?�#��S8>N��i��:i�6�G
:���M֖���nkf]�t9�1<1Ը�?+��9}�Cy]}��IB��R$z��Rs�HP�q�j��WkM�L���1��F�o͕��f-�Dw�����\��ߠF<�_%�Y��s!b� ���Ӻ2G����X��ҋ0��J�/��\U�KN�)ۏ=����XS�|����M��VuΜ��[O���39�_�Hc�T��-g(�'Ĵ�Dv�!B#�7J�7��4�g����bxۼ|Al�r��D�lWzyVXb��訿�Zw_��!�	f
$<C����#3�˸�`n�E�� \<"����8���g|Wg�רXВ���A?G��ԣ�`�>Ҿ�LQ�e�@B�O�.]׽(}Q��W����Cw���}LQl"�p�����vkAo�l�s�2���^��?H�W��i�L�Yl�{l� �7Լy��YD��r��P���xJ��gLԀ���8Ս@[{������w�����gE��n�so颎��9��ex�KhR�2�ߜ���u��r:[���I2GM�B����g������QӐWC����M]&W��v+�t��<5FnӲ (� 
��m�+GrW��~��z�^�r#�cr��<`��(�j��v L�Pc��(+:2��t�V�|c�A����O������N�