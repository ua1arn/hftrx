��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga���<�\��J�ιϛ�;]X1�V�h���G����8(�	<�rĳ 9U�_J���77V'��B����Yr�����Y���A����7�yGR�3�:혾#X�
I��)����+pD�9����������s�JӘ�ǉ��Si=�~w��G�R@���r�m/{SؿaO�H�z%����̐"�>>9U�WQ ������CN]�;ݨJ�diuC��|w�H�-m�0�8�5�@v�!h4��u���;���T){�k�8y`Mʙ��MNM�jĖU�V����A��_����GU{�G-��q{�r��3O�G�OC���.?>�v|A'�6��\�ގ>^�u�I6wj�M�u�LQN�-�ޫjs�ȳ=#.:ߞ��F�oA�N�1�S�	�r�B��h���e{�TM8�o�G���a&`/��L鴦ّ�l����EU�=���7�Ou4��	 ����b=]l<;-RV#`Q]O�O�d�H.�*G�;�hNN�|T ?	m�m���#�&���GT�vMl���[r+�����0���Ub��&031���%���7� ����d]P5�|I
�Ǡw�B_.�8G���ީ�|UO������K�{%e�c �F_M�lZ]x%�2@1��ts�̨cj���ƹ�^��k&5��*&�[[�F2e�t�)� &*��_a���^T��vq*�*3�$'��q�4l@0{*�Z�
�=�xg�f��m��ʩa9��aTNo=IdE�r�Z5��1F�+�8��ȹ�j&/ߔ��O;�j�� 6v�&v�p�u�9d����ܰ�N��(�|��$���&nK(Ɇ]�xs������L�8ϼ,�hߏh��N�ތ�69��"7F5�(E0����v���6�%��C?��G�8V��A:a���@��BQ��|}�����0�ړ��T�, �����҂�j&8��r��C_��xDl,E{�^d7 N�����4G����S|Z�sJ�+S�W�)��<L��e���2%�ttt����6%g͵�"s��G�̧��jM'X�K��[M6li�`_��㼍n�0P�%4?Íyr�`ՑYV�2O����g�`"�J�u]k�H�&'!�Lj�l ���V�4�C�=�h���e,��%4�
�SU��QE���U�� ��A��O,^_�x���y�#�����\��is���9T.Eu e���VL��Fƛb���Ps�5�@���E�؞(@6�EsD��`@T�}�z���A���Mq~�}�%�����_�b+l���C��w�l��S��*}��ӎ�¯	��O�ۚGv�v�:E�FN���G�Q��<9����66S��o]�����M	k�~���&��I�e߬	��C����>��>�K<j�Um�w���D;YL=R��-�����x*p��k�9���f�C\�����Rz�/1����|X8}	҅zK�	���fo� ��P2=G����K��h�ٚ��n�E��W����.� �PsH�-������;JLB�{��x��My��!�����C�.qeP��m���eus��h��f�.П�c�8ƴU��M����-Z�����t��*���}{;(@��1�}��{�1��6�浲ςIګh$%�آ�OA�߭۵�����ӻ�4V�.!*�J��]�s�f���I��ѥ����qNǳ���9�UShwS]y&�N�vG$ۏ��>q��e�Fv�h��Y6!�s�cZ��5�h������!&�Е��E�'�PgI�y�W���9��[[���u�� $������H��)ؙbB�l�[��}tG-����t
�)�С�c(5z���P�4Wɲ)j�N����6�ɲG��<YS��+Q�e��pcD�Řl�:и��^����@ZO�$�f���)Ȉ̆�N�o�Ʈ�>�K*b��*��"�Y,����������*
6ȽIs꣗}:�ı�V��^S`�W�M�����3���k�x�2/�?چ-���)DvɄ:��{�P~�����`sX�dM�(e?Z��B6(-�ǜ�}Q���:�[��xJ���0��-�(��LG>���6
o���֣H��52/��%ܩ|9?3��!6��kp�Cə�_@Kj�_���Α
ˈ�M΁�>�J�1�$�u�"�,���5$�z)?k�Ն�4j꙽q�ĝ�� �N�I�����t�T��vem�1]pBV�a4	l�ν�T��&��tlLT��(����m�q�4�t&g�*^�T�R+��ʲ8 bu��I�y�"��pހ����m�Xh�n��v��A����N����Q6g�S��Ғ6Ŏv�7������#��L��e��D�<5 n�7�Z暐�SV`iqg�\nr���e��j\a��it�̒���d�J� KZ�y�l����Wl�b����V6t��[�J.�y�t��f����Y������E�1�	aa�(b^�NcC�;���^85�9sXXK�!����ysv�E/����UO}QV��*��_�3>>D�.��l����;��w�o7}�\� wY��B��_��L�`�/H� �y7n�J��2]��9j���V���Sfv�4�c���Z��n�zhSr[�7\���r$KQ�6��~�"�k,W����|���P'$�{y�#��5=�>[��O׆�� R>�T�|0�����j���DҌo��j(�_���i*Z@i��'ڭ�[���ʚ�����Gg��D%B�!u$(�i�?��M��u�����ϕX�"���s`��=��Z6Њp���>��ܳFƠ�?���30��O_��4��7Rٕ���K��u����ZQe	�zM�O �s�B�L�B�}��'�^3$�d0]u ��n]��/�>��=X' �M��ֳ���q`�O���LC�iwə�gl�PA$���է&D�,�F
|:�>�1�M5ׄv���.�]ҵ5� W��b���s���PS;��۠�hH����֍���	Z�9�o���Y�ش����=�y 1tvf8D�>�����O
b�K��< ��}`iH�)�	��e[�{����#�7�_��q��� #c�y��ʛ�w�U���$e�怢���GdE����B�q�Y��W���V
�]ҠU��S�~8:zXה��fa���s�8��n�ɼ"�d�;���Y50"��d��J6.%ʉk\v���~��e	 d��_k�x��4�}%�Ɂ�E6��3��f���#���jP�U��r���Ō��A4+zN�X���=j��%�	��qS`X�E���D*/Lrf�-4N2Yf�LP�i!~��L�G��25C��v�j<TW�(�����^nr�?1^a��D�AV'X�|Y�����ˮ�ZU�{�����p��'B!Nj�A��jג��@��ӹ�����>f+����@�
1'.y	�|��o���)�@���s��dt�:�.Y��<CP�/7�9#q�X��h��k�B��Xq�7�QQ�2���C.Eo����z��H�f��4OC�bi��������xԘx�*�t��x!���pu�\�T\颗j"ߤ���䳜爒h�e���Z��3B�b��3Ԫ�H�b��Y���Z^pܠ������ AJ�Rt���V�3/xT�1DK%��TAU�O�8]R��<zv"
L@	uċ̶�֦�q;*ޡ!I��eƲ%a��<~/��F�b"p0�@��k�hj��P(�6��-k!hQ�j�v�"q�/�R]p��܀����U��	s�1���vm>8�}7�
}�đ7�8Y�K�K9 "�`ǢX��"]R�SI�q!�=X&2�>�z&��͖�������|l�R�'~��Ц�"�v�2�~�`A��}H�zO�`}���db��Љ%xl���.€���1'�dw�6x�F�R�,��둤��ٳ��f���>��
XC/)P q\߆�lJ]�c��^�>ؽ�?���C��w��5�X�f)^�e�*���*gK��@<C�
��z�̨���"Q�qjF d��-S����C?t/�b�J��p�[�6�/�eV�\�w�R��u&�̄B;#�<c���k�ؗt��H�z�v§��6f��	G{MT�K�R�� ��)�H_��kP��Yܹ�9[�4���n���/�����=�'^�pN�i����OUԠϗ!J�-=�>�ֽ�ζ����	���tE�D|��M��&�d/���=V���Q�|l�DF��~��{G<(�l3�1J��V86��a\���Gnt=NtvG`�M�b���G}� :�S���O��ԓ�@4��]3;��,�F��B��`X�+�oJ�A��8��ib5�gJ���`/F�m�sU>��\|lFw�5�����)/_)�p�R�Lޕ� ��,�W'�j�M�<_��y
�K��ZnC;�~J������'hqC�>)�(���f,vշ��C3B_p��[n0���$�<������ �MQ� �� PI��2����#ZH�"�޵�
	����	����^`Em1�#��LZ���c��E�߁ڕa�KއcZ���z޵�N#���K.@����a"C�����y�~����o�nz�!&�:��~����X>�UkҶ�l�Y��1�w���6K�!�G�	E����bT�ݕ ��^ &^�9^KD�B}8���sS0o��b��FN"w9�a/�xۺ>�5F
G��lB���6+���k��P��+mAG>���4�$�;ΉW�3S���a�O�+���z͑��XE �D=�p��x���p=�F��@���".9��54�1�����t�귡K2@k�1&�(�HT8'���46�?�k��xu�������0�#��~A]�{��6@�*�x���PT"������z<��7�~X����^�@�~0�g��jj7ݧ^):a�����O����-'8�)��?��ZZ�J�Or�e�?�0IĻ���-���86E}��I]�F��(�4_s�"��s��a�I&�mxQ�(�Kpj0��*_���ѓ���m�BK~�X��}�+u�$��Wc�jy��*�\���+��8\�j�F}"#4u0�f�L7��]%�H*^1���r�샾.�0p�d�3y��|�NA�[!���P�cT^7��V{%�c|���T�W�sԤ��"���r+	���^��T?�C�L�� �h��Qו��y��^��irEP��bH��&�-ԛS��97��LI�d+�KE7/4<|��E�[�)�h�^�Q{p���6@QF�\;��x���k���ۡ�B�����2������]N�zt�� �Li����S$Q_�V:�~��Uc^tYH���xV���R͐a"��R���ɋǴ���@C��4�O�·�~.��F��_�͏���m)��S�sz�#m�iZ9�#kKZTy:oG�5..K��aَ|Aݓ��w�xP19	��I�q@9DJ.���A�n��S5yl�tS���bW�?n��ٍ��H���v��0������a����]��@5䤲�T���,^��8�]J� ��Z�`X��$�Y�l���_v� ��ݮ��������	����O�Y#�ϫ�	̬Z����Le�Zb�����Dy�)�'��#C�#�>oNa{�ט�6�D�q��o�E# ��>.��R��#o���)��G�N]�b=b�::�����y���_[��%�`��b��N3͒��!^��&2�����p����DъZ�3�����7�&h���p֟؈���&�8��&b.��&OW,K�ӝg�q^����VRw����xVN�D  �j�v+hQ�<4H^�om��h����bJ���LxK���B�'E 6y�uT��.��,{D,�n�O'���.���Aw���};�6��u��#tD���&��tb�h\���k���.՟�ȳB����ceyme4�ɞޢQL�ܼ8�ˬ��W�� ��UX����a�YC�Λo�+��W�8����X�Vq�ߞ@2+М:����`����㈣�	K��I��p�H.���d&% � �0�tagL9-CG�<�᷈�O�U�Kɳ(�	uJq��I�?�%)��U4�y�%����B�@Y �l,�Y���,���F5o[�׭��5ٌTko�����0�2��9-�mϦ��X^y�߲���oH*�D����<MV�K��l��o_�x����c1�{��3�)L�|�����,���4� �(�R)�$�/�{x�����y�7Ɠ��9of��G�y!h��.|�w��y8���.��n~��#b']�8r#�R���Q��i��	��Y��ݤYh8Z�n��t��<.O?��j;�f|����������p���E����ަ�Ȣ
�W
����L�{�	�u�A�6�������(�䨫�6�����������;�@�Z�dY��Jc	ǭ���q�&uF�9��ڝ7R@-MyS�w^m`�6������n�}�K�G�
d4���R�����w6ZD<����v/���\���d�v��զbp�u{�=��/L#k�P
B�vOX��O�v�^���>� ���N68�z�_Hc/����۽����#B�I[`,����!��$h�f}!�P����Ie` ~E`��!�����A%�
Z�*�����ྗ��|��d�M����б�̵���o�sJ�>T���A��T�^	K����{_ԟ	>~��9�ãsx]��a6�����˛Ȳ��D^ܥ��2e��+m/!���sq��0+�����b���\�5���WV�n�ۊ�x��-F�=�4���k�˩Q�f��)lo ��H�t�G������ ��A���o��e"� �����(a�0�00�q_���vcY�E������152�(� S�\���%��H���6�V{�ܤ��+ǥ`�F�A�u��D�b\�hof�Ŀ5"�&`�A�^o�DC��=a}�JᝇrۅS�yz����L���2yߋk�C�cy��E��E.��W���7�A�tՀ�M��6���꒒�Z���W�YJ>#AGg�U���g�y5�p��H���,|Vd�@ ���c�tv̢[,�{�5�o�w��:O��*�M9�$�2{�Taqcê�����6J�[�QЮ9u������ӈ�57a�v_nX������ �ݻ}��J��Y������R�
�]���,���� ��'C��h1ᡡ����sz�BQ���t>f܈��kk�Ǜ(zlɉ<��@��i<��9-z���2{�"9���M$���-��,�3P�ߎXt����P��� �Y窳n!�|tu�x���~�t���o���5軺8U�c��`��s�*��h��^�Ȩd*"G����*��:k�k�e�u�Yݦxx\{#�kxpL5g�l��U˪�^Ie䦏<y% �HdT)O��O�۽��p�(q�,6O�ޣw�_@;��M�}q��tJ���ji|tc��ϕGw�R�"�X�	D���xy����}�N$�(w�ƽ�Wt>L�2P�HsB��(^_�7`�s[?�L�V��n�z��o8���B�
gb�6n�r�,����̶1�w[�gTn'eىm���|���.I�� �\�>iy��A�[��e	��:��w»�$�4$�00͛4�C%w��ۉ�4 ��(�v��ĥ�0�B/��2�T��f�\>oν���|pr��(D�j� DO\<J��"�*����4,��	wԿ�
-U�_��^HQ���aCx A6�,�/K�[���F"�³W�(�۴>>���V,I���V=ǭqu���6�t!F�xKC���K�f�7��M 0..��}D���7$2*
�h��a�����������Q�xs���0���U$����7L4��M�>S���d��AF.����(�����ؤ��`j���eA�T�%ZnEjH�^�[�zQ$��� ���HwK�(���la�mه7����+Eˡ��ZeM �8b͑P4:d�5��4�h{�8�%�J��~����Ԩ����=�Rߑ��2����n�F>lF_�����	�v`�[��^(�%���KI0tJ\��U+uqz�B-b� �IJ"¼�p���+��:�J�^�ń��ɑF-3����q�?��AF��0"�r���>�񫔡�;4|����6!n�`
G�ع>���Z��+��طA>�1۾988���l��c閗A36��)v�-�_��hmHZ��5z?��˝�O��i�<�2����෸�;�-E}����Na�%W����=�%��� {EFEYa��0���:n�㼪7H���iBqߋ�+D���(���c�ݧ�]\Yszj CbG�0{�J����v)�=/�G��Tn���h�*M&�h�'z ��n���zo����U�h99:K���/���y�iU���"@ө!�m�Gh�|{:&��+5U�}����H�x��` �ҲN�P�D7�W�{�ᤀ2�Ki�T�)� ��ܗ��ܦ��z��W��C��D��Ъ� �=tΣ�1��q��Fj~�a9u�*�����f��g�	q U�_w={��wzCk-�^;�n�\m"e��K H�k�����&���\׀N��8_|��؛}LZ���R[��v7~a������ձL�>Xwf=���!�O����1�Z����`�O	7��`b�6��h����Z�A����� ��;���c������q�"Q��+�\W!�B�m����۲�����
�3��\��.��뀊Ƚ���@�x�5EC���;�Y����|���\0����D���c&Zi1r�Rȧ� nΪt�d�����t_[�����5�?�U�4�]����&���Y-�RB�� 5��ʌ¼R8}/��&Q�:�~���<C�vZT�|b�ݪ( �.�ޮSMf�T�X{�G�Q3�����f;�[�3�Zo��7�~��}��W��И��M�c��q��qd|�qd�
�����T��!Л��k�n^��ߙ,I�do��Ng����G���m��xĈ��fD�bAS�s�N{o��Z(��mi���d��(�>Oi(̙WN\\\8I��H�2��
Ts�C�l��>�4��1>bd5.X��׍Gm��
:uy5�0�s�ï}��l>�8���z����'9e?��<��A���Y�''�8$����i2�
S�Pd<�X��xBd�<M��,��7�
��6��O���|�A2w2�~$)��
`攗mt��G�5�<࣢g#���HPԗ��8�D� �.�~{��\�*�!kg�h
�rVƞ��KL��=!x	��S�J�m��4���H��BY�6��ۡYo�RƠI�����Zױ֐tpd�f�CG�_��60[�/�-�8P�y���Ʋy/o����U���h�@�C$Ǚ��i��qߟ���m�}3j!��!�g�\��DA�$\�����J@S]�ɆD����-�@���'���*�d'�Z�� ���3I8�Zl����Hd�ε�x´ƿ��`@?ʧh�U"ϑ^`zW���L'��ũ�W���0�p�O�?����>f!��Oӥ���r_��{���`Ʃ�Y���7���"a���W#�+-e~��6�a��观�#�8,��o��Q��1֚K{�cR ���\n\ B�i">�P+2Pr�,'$��əB28F-K�w�P랃�{����^:Į��b[t��t҅�v�ί\��0R�H��Yjz;�1>K�T��7����<��b|��Q�;j���E���8@7c�,���b@ȫ�!V�aKR&���F���-念�Ac|���9&�����R��MQ~�taC�,�%��k�}�Ee'�Ԁ�����E*��B�y���<Z��S!���I�Nl���o��*,��0�A��h��.v[��c��؉���T=k��`q�t�T1K�.ui�`�d0�T�3��k43U^r��M�#f���4�?�o\Y&��Ü��}Dz��ĉN�9r�@�#wր��������<���H��:�������,]��JQ-<ް�J�0u��� ^N���hԁ{�׆��H�YY\�����b���	��Ǣ@v��Z��O�/��X�P���/C��&U �� ������!�d�mV$�����s�s�������z8�V6s��ݩq*q����L0f�������a�ԭf�b������2�lG�v��\��RJ�,Ɠ��ě+FXn�`�d�N� �N�Z9�9c�(ɀ;R�/��u�Q�~) ��k3I�ʝk͆+����^�<eWQ�eتfm�s��{��-��%���cp8�Ec��⩘���ܧ":y�`nx$�;���kh����/E4�ڠ�6D#� �m�3u����h^�:¥����Y0ר.��T,��{����R@q'��^��b���z�&�(.	��Ie�"�"���_T�ӏ��9�"�	���F%�����_v����g�������vl�/��U�ĭ%/�ƧnqEd�,���8v}��I>Iܚ�n����� �1����Jh�"�c$~9�M��C�Vc4�
e����R,���3�[���,��i�G����@�{B�P�~	,�o���Ԕm��7l��!�J��8�.���v?�3m��Đ�,iZ�dv!%���m��;�j������gq[5~�[�\�F����G�j������6�Ld�m5%�>ZT��0��)��
q�=d�iɝ�_���ϽO).e5��p���5���n��/Z��vֿ�-�qm�S_���ftd�	��UlXτ��T��x�D�/��;����M��y���ɬ�7��Z8�cg<�Ω�\�gB���>s��-�9@ͩ�j�D\�x����J�E�����x0)� �{�-���v��X�;���V�,�;��O�"Ǩ}�E
�y�!&H[F��r��p.�>�AXI�l���S�]�MfN/lk��=y��Z��Z2�R�_h\�`�%i�@�e_�!���T,��Ë�/�ɹ�*�}l�b�$�'�mW*;��F��T�� ��m�='�K�q��<�����B���0IZ�hŅ�K���Daj���RD�W�]p2�K�Čv�洃��锁�ً�b�`�A��S�n'T2cL�2�`A,�dOmr}������y������IN&�2?g�n]�:���/֒��N���._2�������:54d��<} ����5qĳ9�d$hО�U�ĭh$����	ٸ	���@�:��|'�#��������ĻM�;Ã���Vb��r0�g�Nm��^0=-A������el�ᆒ�zUo���J�$��oE����Wi�����U㭀�wG�r~��<���o�wm�e�ݳ%��'Mb���v��22u>�U�Z;�˵�i~rTS'-�kK��*ꡉ`Z����I� ʂ;�`�v�����g�'�w��",i'�Sr8��*�߰�aӚ�?���2@���v�!�׏/Y�t���.��o�it��3�����Ѯu�:1�""R����R�*���2�_�*[�K9�7���s���x��� �D�A���䙮4�ߚ<6��_�h�-͗O��D�{x���h��<��P�uy��;>-b�����3�6�E_�#��R�`i��QcQDE�����Ԙ;��6�)�;b��{�|�n5p�5sOT[t���Q��S���d�p��4��)?}������@u����#\M�LfӠ[���gO;��S&��5%�Ѧۈ�wpY���)0�ܑ��r��'��H/�T���_J5SA���D��yiL��]�i}%7�/ߍ-��̜n>.h:������u�r�����Ē�+�N�p�S������-��T�VgY|��W��b��=ll0vc4�]XO-EW�d��ns�R[߽ݸ3��%榬�̗._�z�`��FO���e��{�x)C�!c;�����K�A���]�P�E���d��_���:��ʡ&��������	��`6æժ�/n�T�=��t*X&{}U�B1��o�u��^8f �΍�"�+ǐ�wxw��w���f��h��Y��>g@�E~';�M���K�sk�јU���,��C�)�Ё����$ދjOS c������?�"�h]X�����%,��)Y��=F�W�<�T�4K��,���}�{��@�\ �eZ��Bm��aF1�Jt��M�Y���l�'�it�;Q��u)n������������k�Ҋe��?�+�Ԝ�g� �0���&�Ս^CjښD��-��p�<]tֶtŢ_�b?]%w�\b�����(H�sa�a �0���n��݄�UYfyX1��-><���z��T!gC���K�p�"zš��.�����~iM_���)��������$��$��eE�}���ݪ�ʾ�w� �e�zh�oe򯔷��8>l�5%�b5�t�Ho�)/?��rS�n�
��C��Z��
���:>�"��o�4<��z��Ψ�2&;�4Ƀ(9G�ƙ��%�W���RO��_YȲ���lT���ip�*���"?N
�9Q�ά�,mp�($�^�e�É���ўx\�g>�%��0�;a{� la�=#=_k��l|�cn>	_�H��UB �����(�lY�����F�(!l(&�5ݖմ��+F���|�{��l�2�r�v��{M;u���w�|{�.Ip��_Anb���ų��#���@�B�5��uj�,���һ<]��Q�W�ah�s�<٢�鯪$ p'ӧ�gpk[g�G]�q�� �l2\r�:�!�j��7�{ϴ �!Ė�6�@xC0�#� �{2}�X:�E��˞�:��37��ci'>e��,�n�ada�S=�s�1�ێ�������C�͵�岆`�n�h���۶� ��xyI#����q6��!bL�|�$�)���R��n�#����VJ��0� ���q@���� I��0I�j���-Q/p���n���ؤ�� �)��	|:�9fEy_M}��o�Z놶1��w�j9�<����B�/{ �}-#�d�઻�<�u}���z@Z���5��}���$I�<ӭ���vnU����p���:4�Q	N	���]Q{�DTɣ�P�l��g��y$DT�����CZ�k c�Z����0.�{�AM1n��������)���6_���u J�!x���-��m]f�jM-.�j�)�OB6�v)�\�]�3���Wy�8\+~a�^�F��e�M#�f�2<��ǝ��w���N�-|е�_튐��Lp��	[S�#�`�T#QGU���&*�����.�@�[�x"�D�V���V�m'�E �:q�K����6�r�8��ʮ���8ɳ����X]m���;�X�8�)��^G��9s����q��{���it�FP��ʪ���FF:�씳o\)�3��@�@^+!e�����	��	@kD0��<܁�Z���Uڷo�7V�`2�*>�_�s��R��B@���_�b���N��ɭ�hj��WxK6��k�x$Hݗ_Ż(4���&������8e2��Si����]���>_�ԔTC9\vTr�l��'�$�BPY���탣�����"��{i�s��
��t�����a��!AH�ۗ�)g��L�ǝ�&-�kl���Hd�\���W������P%ut��|����j��[W�=	�1>�*<���9��ʷT�x���n����sH\1]O����$��ӑ�o��f/����'�+׫���'kW�z�]\�d����D����<�����Ð�Dp��e!��Ɓ~"Q�ozy��CjA!����jtFD���[��M��V��n���Ͼ����� h��Q�ߐ�/Y��8���������Y)F�f�ece�������<��bM�u*��<[k�n`V���|���c�x��h�~��V��}a��d��O�ċj�RF�d��/�9����eN@��<탨�@݆�L�:u����c�M�lM�[LR+��2�f��am,߼�)A>Zu:7�\��������#���[p�s
Z�V����yԈeQ	�nۅ]�y���=��K2)�G��X﵌�%r��Y��	��!��ӻ�L0w�wހ������Y(~�������?�x��iKrˆ�3�_��E��|+��"�b͸��=�cŊ��y`�~25}п�yП��1w�'�[�E]�,xv��m�R�%7,e��Y�T��Ӌ�E��� ����'�"�@������x��!`�����M��hy���+_�h�w�-��o.�6���DD�fA��!m�G4"��T�9V~�/����,�7q�
��z��֛=F�W�y�Zy���@$�G�q�^sO�C�m��p�e�}�aD��d�R�� "Ӵ����D��_�a))�:o_!!3mX��lCT��O]3nK�%��3�@�����7~i����.�KL\����D";G�G?t4�5F��*	�Kf0�"�Ꮷ��g��O�18��Νn��wIw?�)؟z��n��ozEEd/����L�V5"�5���ř�;`�O�p��)�����6W��������&x���u��s��RP��O�D�+G�z�:�CiD��f"s��m~���P��q��Pң�0��6��.J(8�1�$��j�|Z��RNV���f��np�y֚4�Hm��ٸ�e�|�
�E1�B;��B,ʩZ����(�	����9#������%o�;mNZ�[��F��_�~D�D`�ވ�<5'$��s�fW���.d˙�>�	,��`g
�6lsջ-^����g�E��x���5����U��T|�m��K�i�wV���_O/��.g�������������L>��×;�ZS~ez���6�i�����ն�vB2��H��2��;c~MX;9�ԝ�����;�FT�˴=�a�*L�L����.( ��m�h��PT�Qyam��d��2n��0�Ѵ�:�y�"#����w�\F2�� ����&�_�ɡ�;@�l\�:`
�x��햛������d���i�	a��:~����C0*���.��6�
�y��-��5T�86��)���@��J���@k�h��_�&���L���BPBD����6�,��S��<a�9A}�mvD�/NSyeu.���7~p��k���LU>I����˾�]�B�E�n"|p��x��^��Q�YS�Y�8L�B�C�x�{�i��P���3FB��y������
�=�;���t�MBÕNmdL��q^�/UM�;��,V��ܴ|�C��5�p��1M���s�M/��W9<�O�K���2ˀ�����(�V6�������$+&;(�:�����U��;Ps��*�`Y� �=�١�OM�D�����K������]���"�6��@���S>��?������k4A�l>�ڠ��=�=��V�Qo�Ό��@F��Ťv] 1��8�)3��뺨 r�(�דk�"�,�m2��m��wK��-�[E�/0}��W��R���|�f�g�0ɐKo\*����N5_߱S���xᓺ��N$x�I����2�ϡ:X�
���,�ن�E(�.03�@AB��]�L����aՒ�g�SP����[)vM{PP\	j�@p������|�n�!�@wJVf�W�B���8z	(�2Ȳ�k/�΍aZ5/���1[�:v�$5�S���(L�:!tB�ct�ݦ��:��p��ć(a�2sRڭ ��t��gh��$��W>�n����5V�8�����v�8��]�p�Ꝫ�ح0%b�+1��ܠ�(۠B���;S�ϡ�e��ې�暊�Y(���� c|�d)�_�����يG//�\,�6���,��+�h?z����:�Ygz�I]�ז��+����A��6���c�Oy����=qՕ��	��,d�t��v��9�/	��"\86>��9�Ꮾ�oǜ��Œڛ`�Q&��:���Rr� >�7E۷�Gy�tR�(��H몏Ht�E�ո���ڤN�y�>I�:!
,MMxB=׺w�������`G������m+I;���w�i��Z�_}�9>)�{�w=ϴ��� ,��2�vF���~p{�yJ�!! z#�4G�G�ҬE�M.><��e�畃��2���}NɢB�w�fݞ�E�iQ�� ���`q;�eK���֮j�9��-��/\�W�_`�8X9��H�,�xNo�( =X�3�4R�q�B����V$-��//��=��2�ߡ���ݟDQ��6-&%�c����}sD���pY���d�LP�}��`�~�Ho���1�c2A�����3�&kXH�;���ʐ@#����Ȼ�A��MH��G�NÛYҹ�E�X� ��j�NS�4aS2�XB]K�����(�)����QM �@��2Ym/J�*M�)��}s4��N3Z�1��J�lE�ɪ)W�#�f�]��0��:��!�t]�& -��[m�KP��F�J{4©va�؄�����\�xη����d٪�){eV�K� b����\cZ=��lu�<���y�_��1��`���复	*
�l%�Wl+���G�lh.���?�z�D�#����<J]N\B*�?�p!L���FH8�g�NRN�T�{)p1����>!f� f��)�;Y�����?��+����U?gD�]��q�Rxk�[��z����|r3(�!cY�,�e>����<5D��iG^�R���UOeVۛ�N,�{DR0�`>��0VX�o�m^���n�D�0�����-���/����� p��ti�=��E,�N��nbE�T�Vt���ȟ8M�3Qv1_���BBY6D`.��W4�Vˁr����$ٸa���ha;�xiU���ve����'����.�<�r_ V
P�Q����nA��ft�/� ���#z^
�So�����s�R��,�
��)�D��p���3@}���1A����9CIiXvO*�Δ�6�y?��}�g
�o���a�Y\�_�^0w�چ����i�s�:�����޷Ѣ[eq��k���
�2��~�Eh��;V���f���b	����G�f¦�A��=�W&N�hПq�U|�*çw��a��P��|c�~������A�n��̧�;+I��s?����ABr�+�饇���v�����,�P�������@5{%T�Ռ��GBi��){9���ޚhU��Us���?�1F)WApY���	��D@��W8�l�;�(����yf2٫�5��zh>xE(M���H�E�s,:f�ﳕ���3t�t�MH\e��>��HY�ɸ(�qT�Ve��z�V�˧�ʣ�{P�t��Y'��^V�Y'����x��X�_x�pM�q�V��Y�ݻ�KVzk0iC>�b��ZL�O���ѧ���Q	��xv9d���p�m �_�Ye.\J��|���D����&"iWPOzƔ�Ni$`*�½���z=�O�f��8(~(W>�p�P��`�vq+%���qE(���� �=���
?���@J�tX������:����n��&�`׭�~�g]�#��RP4=U�
��y`���M],v2ec����ДH%Y"7븑@�;�����ydX�Nulm�;�!�f��	6:��8��ʁH���	q @�#E�PL|@�pVp���r{�h���=�'�Ko�pma�(�vY͞	��8���w	
j��j�+f,�0:�b�ė(�O��HH{�a�$�6E@��i`����:="���%L����s#D��Ks��ж�����t�HS�L'�\;b��XzBH�����9�KC�^0��D[�fS�ߍ�F�x��Oܳ7 D"r9 &ɂQ�8�YL#�jޠ�/Ƴ�3�k,��9q��p�#檈������*��!d�?�,z�Z����݇��T2��:�A�h�Q��%�9�b�;������Z~�@ �����)�p7�۝nfl2�fX�ƕ����ajt9�쪚��q���Ā���g��b{�8��\u ���9~�'ߣ%����~�ղ�<�F����i(JOz�q��L�:�Mı:^R���T)�bh-}�+P���D/ I�>�c��m�/�U���+[9W(�0�i�}����}��%~�u ƿPeP@'m�$%��i���0�v"�\B��qs(�6V���v���:h���+)��9��	Q1
��pxc�p�بq���R���J�ѥx��e#�{�	�R�#�8�@ǚU�0o%f��S�CɛmǆT&�������{.I�kM
�/_��1�7��M �l�c<}�}n�/��Yךl��v6j�F��*D}/��ٶ��Z�@�B[/몎�j��E���[?|P�Yʱ�^f>�eI�����z���: ��zC�P�S��u��)q<�K8�Μ�D��dY!���$���Ȣǉ�i�1�f��a�\�BO�E��3�J�WPǳ+ل����#S�O�2�+�׫Z@F�_�����-�@�%Rr�O��՟\�U�/x;��@��g����J{��A�^e餂"3��X_��5�(�l��z�.S|���E�����MF��r�i��*�JM�������7T���c�/��1_���'��<��q݊�²Q���uJ���;	���*�<��'t*���(p�3�qs���4�C㸙��s
!I�
��P�<Hא���� �-��1�7�t�X6\��2I\����U*Τ	�F�{ڸ����s��������fТ�,���"Ap=�	XlBj.[��o�R�`�$�!�%	��'B���9��m��廓�F"S_\�F|OK~����[�ڪ��r sy���a�R�������s�R��{���'���^�6��c�O��`���w��P*�Q33����eoƒP��x���ʦ'R! �j
� ��(�E�Ju.o�3)��+�N�t%ٕ�=�D���3������vv�cpuǮ�!ޕ�]���ª�b�Y����3V�C�Y�����l	A!�1���I�YC����p���*�aQ���L�i�q��"�2�Fa��xѧ.�a��y�ts57e�ҹ?�b���(-���J�_-���Î���A�����|_6�:�/bو�$�g_e�햷�����_��G��J��+�|XT~$��LkG�B�i�]4k&�&�s�A�&ᱪNA�J���~�ΰ%�T��$o���<w}&~5ne��t���ѷ���߶�練����C*��D%lN��;Y�,=m�a;�k�� Q/i��~�\C�����O��(D [���F��q`}?�	�j���s�$�W�@]��MM\�c���d�����B��vǲ��#ťӌ�6v� ���}����)]�{t�=��W'�����̊ױs�T�Y��{�v���k=JC��G�|�Ba�>��q�f�|=�,֍���*���V�ڼH������d��Q�&ُp�g/>�DWDǊaNF�~�ȸ����������?�d��T��o���ʆ� ��A/�E��&�+#<�b񛚋-`�ڐ��#H�|�	(!���}�� |zg�[��'V��������N��Y1I�@��w0C@{�܀���?z�����{�Pjt��v^t��8�p�|���+{ċ�t��F�ai���8��E+%
��kVm�:R�8�k��G8F͏O>(�����G��dѭ7]�
��j	�I�2��]7���qTϋ����� z�hh���~Y�i6;;ɟjҭ?ܙ�Hd��s�BY�qI��V��6������8Z��n���iUU��1L���k�p.B�5g�Xzǲ�$��0��4Y>\$šK%Hd�z�0�E!��'���TU)9.����ހ�;���b�29L(���46��BE�%�"�mGI��;�V:� 8@ph�c!��_���ʜ���(��B��x�bD�W��K}�������1E�:��{G�+U;/�I�ż��c|�i�^�Q���k����6-���~�D>��bh)zw���V1l8�φ�O:��:��IL3s������V��z&�߶$�9Rcj1�ד�U�|�v|�K9��� ��f!>�(��s�Q�7!��h�c��<Qv�X_�y�:�XZ}׍�Cd��B��t�cCf�MIh��Z�wZ"�sSV�S?�BK64%���mtg��L�v)���UMH���n�u� �d:��;��"}�?['j���'�v%��[k����A���%��cMӨ�EKb���	��l�-؆z��D��[ %$��Ӊ�L�s|�-'�_�cQe�����v'��q�ҕ�=}���H��{T��-S!S�&��בa6�z4�^��/1�#�۸K�abf����[Bײ2PV'̱O��s�i�U%$Z��#�Fq<S��qِ��x֊ݮ�<�iw��o@�S��5��S�NH�/4�%E�H?�}Z��W-,��v��=N�G���^�~x�.z�O��u����_��dqJ�I{y!�x��6��V�^�ݧ��T��!Oֲ��� u,��	)���̄��*�A��35���E�W	�A&�(�viv�MU0雤�nx �7T��B2�>߀Lv@�ޘkj,kd׵U�����mh�`#���7�]020<2x���5��׷�Λj�2%���	)�9#�������Zv,�zY�Q���T�vZ=��#MQsW��l�V���1J�Q����c-�N�h�J�.+p g��?:�g��L��ܨ�b�ҖW<}֑�����r�;�ZV� 	��a�9���f*@��j����eh$ř���6B��G��N�k�^sā�@�����}J�/V�w�9���r	�>I̧7�[H����ą��T�.������@A0�((.a���%�fc}-�h6``L�}�P�G���N���E�l6'�i6rA���R-|x3o��+��,N�,P�z �� ���\;����KT�Ȑ"���7�/t_2ci�Wԍ�w�0��1&j�6Lf+j[��}p�Qhׂ��>XqI��W���c�!��qPt)��8�_���@�H�X��G��66S�qT��!�2���r�SQ�(�8�#r��#&&2�.Gr�K0=EɄ�̣z��I$2�3N�>�����WI�}�^�CGm��{�X�(@���њ`9:��9>��ũi@�Z����w���hԦ�A��np���@TeN�_SH�FR��o"�`���
�\�N��DP;�ڄ����~�?w��� ⣠ٯ2�5���A��!R�\��<6�;V�7Xo�'7��L�xʣ��6��c�В��8] �8���ח��% ���)�L�Z�����:e-93��$R�>CȾ�_�!��F�'�v��R��N[��>��%���w��9���PAN"Zs�|o�+1�⫚�i{���q+:��8�~@��Q��]�պ�����я̆�  O���vW�҉�-6p��y�+OWU��I�9
_���xz�|ͦ�G{�8��yo9����R�z��&i�_�+[V^�+A����1�P���t�f�.' @DS�*}�����M��U�:6Jb�������Ģ�����	�.rV<�`/��;,T�3��/y\��f�a	1w�K�������'�Mɩ�T1�S���F&n���?�{�އ]g�e��4��&8��>�͜�~b�gRK��.С�*VV��s�+���NM�g)s��� `�G�:�W�x�s��r6A1M]X�HF��7��:��*'9�=d��<���둬����\L���T�4K'�!i�h֕�s��[��C[�|�)c�qV`��FR�ϛM�ժ�O��B��,���65@!����Y���(�������Ye����7��@u��p3��9�GΏi��z��$�=����a2�{�yT��� �z))]D-�BP�#�wX�,�h&T�mO�Z��?�I�1��,l[8[[%�z>7B��øb���L��� �q2��`+��꜄���[~�/�WCyUZ�.T��l�-�wPp��8f�,��G���J� Ma��垀��b�u#b~%���n�:�P�*n���':���#4��
(}�!&M@]�A�&>�I��.ڊ�B�hUB��#��A�ހ�9KW� _M֡�q���r�~��*�%�J���J]"W���~�"�����	K�L�זi�����R,}+q�}\�(v����L͛��;J�h/+c��YV*����zK�j��b𨯕���)7�`�4��"����:*�&�?U��a����x�_fZ-S�bRs��Q��ڰ��'��]�JJ!�ݴ��yK�i}o�n���Wz��r'���NF{I�'��-�Ϊs�Kż�Eq�(&�ӎ�9���s��Q��
~�{vr#Sk���MB�cf�B�/����ưB�J��̏�������ݐ���Q�=]�������MdjlÃ�Dw��0�����?���n#��,��	����x�!]�?����Ϣ���r��_p�p�:�a�h�s���J��W�����!:�q�s�ЌX<򫠴�źW��!O0a��Kk�|鄤M?���Ȫ�E����!8W��	��k��o�Z�Y	jJ{?OK��5�Ѷ��e�D���3Aϭ���1�:�8p���-0c�5��c��
&���\��rH�����|�̣E���h�^:�w�s�)|���ҁw@�v �q�����7�"��X��h>�� �ғ������F��������hê`ٲ�b>1�9��c�UG�b!Xrz����"H����	#b���\���'A�vlבŎ�}���޽�fɕ��/����`��CRc�un�I6qi#�O�ZK������t�C���s�=/[����Y��.ک˺-�;�6h;��E���KW ����R��[�J�%���y�2����ERSHHG��idGu�&��L�D��#a�RI�k�pH�@.(� Ǳ&S��&�jŔi)�$\�@���28�s��֫� #�"9K�f�zSٿ�*ۙ��Dİ|�X\��[F��U7��Z-�^�>8,�.��j�Ո��M��Z�n�J`0��p_��'+�Gd-#����M[�q�/ѾW�!�Ӽ������9p��/�5l�s�DO:��yҒ/�fX�yF^���-V�A�~�Q��\Xk*�J�����d���]evӹ�#��f�ZE��+BLx�@GnYaw��m�B�$f�yJ�7Ȅ����k�W��=�T�kY	P�騇�A�
�`�h�#�g�Ɏ����uO:v0�E�]�-�΋��<��^�+��K��2/��@��D���_�/�/���Ք�����O1�����ü�ⶁHy�M��j߀2m3\b۵]o8Ν	��O��[=�(!�ӣ|�d�R���9_�.�L��C?P��4�Z�f,�M!K�������=�UH��L�FZd��J�$��a��<�3t�S�:��?t��GWZt��D�L�Vg�,f:d@P�Y����=�h�����)9؂v"eAd"Q������xH+ϑJeI5Y� nF)�y3�+�/�s�<�_I�<p%�˒�����$Ȟ�*Y:(1��U=G���M_֟��x�k��gKH�[[e(q����/�p����$A��¥72M(	�xg>=�.]F�g� Ib7�I$�K�d�[�R�L<r�� �����F_5F��5D005�	 #���hVj���,t�r���-H�ͥ{|��-��M��n�u���%m��D�o!8���*���x�+�����m��H�`�V^�w�wJ���Z6�	�:V���"a��a�u�[���]��1E�%�k8A��Ը9�߬b�gn�4ꒃ�lTEی�_`�9g�j�C>G�<�_��q^ �j�}��4���S�8�E���h���l�5���]ŹsJ�6*�e�%��Ld���/��t�>��`���"$�3�+�<5i��X�.�rYx���LE@�gp;pyW�������h6*�EOfA�@�����W��l�"�#k��`
x�縓oc���K��b��E�����Q�95.���3������������8�K��L�A�?E{�uaw�O�n�EZ�=qK ��:q�Q�g=�t����!I�
�8��8�&��^����K�1��L�rיY*D��1	S���HR����\����"�S�x4��f�������5��y������G�����e�Ca�\�5Op��ϿXZ��^u:����
��b�����$t)m�� Zv�'�m/��ږ_?J���{�
 ���,# �����=ds�2m�<F�-�ĵ��~�e䏄��}`��D�固'�ݴ �?�����QR�|���L9OQ�>�6; -��Z��m	p4��Z��[�&���D��F恔}^{�
u��bT�Y�����L�ќ�Yw���{�����"�w1��[�@?�F��\�]�u'}���~���z��J8��`�/7�2<����}��{���V����-x���=�X��wC�r�X;9���{~�54>�b����i	���8��p��:AU�����f�'=�+y�e��mŅK#�u�Q,�c`>C��#%����}F�-�+[��3cA�ß�7C��kxp��/�����&�'��b?�\������#�_����U�X�R�q��Y�p�E�2�f��#�H�X��V�5�%Cx�Il�	䨾Ia�	�$�E�-�O*�W`n}�V�m`��������TN���HO=I:���y��γs��B�o�?j05��}��Q�UEP��}kJU_l+��&�&�0@"U��p���d�"5���V������3�y��b{���ۘT���T�>G-��Z��X�u��w���b�%U�w���{*Ƹd���*�`�g�v�o��ŕ��Tb���u�Kϲ�f��Mt)su�U��6�U.Ԭ��p�!�.jP޵ Y�B|�f	�C���1�X����Kj}C���e�.�?�Q-Lb́����UTպ�Ѣ.���TbB��ϑ�����ܡ�.�����1�o�D�mu�u��HW)����t���̥+����nH�,c:%Q���P�4ȋ[[�/B�B��v?N����F��6(��d
!�A.D�u�Ȓ�Jw�Y��/O�<�Q̎��8�8G��Jw��ڬ�w���̙���~�,$� �~�> +��FH>\��L�H��N��4�h'�����dNx��c���y�+�Ic��(�rb�t\UE7i��-�tW-A<�^�l�C�%f��=�^`�F�9FKe{�Z�0�Pd�����Z$I�F�� O|0�xi[�>0�K��w�ab;'��\����=�`%�80���}�^�N�Jcm���
���[�Ԡb&Ȁ�K