��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d���O�2 ���b��$%m�~�Tg�(zx��{��b�C�M�*Y���9�<�,ҜE���xKW��*1��	�]��Q���Lt��״E���鄇)���Mv}�ch�E��]P�59� �dl��� ��l���dm��Q��)�1��e�^���ϕ��Q�AZ~յS�6�4��?�	R�9J�s������Vٴ|k����|�����uz�Q��H+��ezh��߲���1Y�@�;�5���LȄYfi<��c]ʬR�e��n5I�R���3������D��%4V&�N���GN��$=o-�AS��4xD@���0��{k�����U�B~��j�K>v����g�ɢ�x�M/<�L��}*w@���eN=��l�|T��ܒ^z0>Z����t#"H���V��LB{�$��߿o?!.�>-�:u��|y��~�� �;+��ӌ��&�g\K���O#SX�4�2z҃7ӶبݱQ�U��PD��h�_�J�ka�̐�;�a1k6�V�)�A���_�"e��[zs��[^�2���4NF�Od�|�̪��p-�u6W::�Wsֹ��Ԧ����(�ș
�j��` L����>���b���{mђ!N��t���!=*|r�D�z��g)�5��K�^ �mm:1}H�����f&��\�1}�4N�h��,b��D�b����B�{�S�Ņz3q���G����`� !"���Y�2a�'��.�����I���g���?*x�H�6��Ǽc�nR��6���f<����v���PhX|�p�,k�)���r���&,.��JOi��]�m�/�K���2����2`��J�i.�'���֤�1
���r�_�;������摐+�����߆L����Iu&l���@d�3x�i���O&"�e��쉘�^bvAKƐK���8��Χ��AK0Ü�G[�u�7��lƒk~�1-0 ���h�;&Zd K��`u�B��:��Ru��_��;���U=�[�SzY�a�j�ƨ+�ܒw	بv���b�rxkiVG���X�J�yy����2�c���{5宀�<B)���5�#pO�ǻw	�LW�RP�Zt>��!��g}�Ϡ��E���n�k쮵L~�����4ʊ�`�( ��@��c�n�<���!�흝�g�A�;�۵/F�Yǂ-������hc5y����
�-��'�N�����%?e&8��P�^R/dO��3.SlI:z�e�l��"[@�PZf�3�����f9V���"���=�Lö�ܭ�;��8"+	7V4��Rę��]�|:w��
8/���8y�Ҟ疸�%H�w٭	[������-x��0+�.B���W����;�-�Y���z��s�Zҍ�M���t�xu��^o�Uh�ݐ��'�T��U�G񴥂��R�m,J���}8��x���������j^�j���3c������z����(h�:t�\�{a��4�5�;(�#���,ul̆��'^�$l]����3��
�أ���:.C��ȵ�G�o���c�@�J���S`��Mt����(>(n�W�M*��-1�u�uU� ���@�qK��<��$Õ2'9N�j� �˓�Oތ��ddè!�J�
t���F���j��D���������ͭ���������X)���"�w�`��1��Q�x�-Т�L;ɂ'�S�{��Nx���x�yR��z,S���)j���JxhR5�&�\w��U�ȸe�@��ߌe^�x��gf�=0-���M�̻�@�h�8�\·�o�.Z�P�/�	Ν؝^#��"!9���Pxf�Ȭ\>���,'&�7���s\���;�\AIUE.	[����&������6 0�i7�}3f�8�����qdI�?�Ai)e���r�{�	����E'XNݗۉ�DJU|������I�$�6NEl�N{*?R�a��m��5�@��� d�Io ����p#"��}�|��;>%b���,�B��^�d��q[���3�wvk�i��A�єY�c����N\W��kr���>���3
{�4d��O_�%�oȁ��Q��w]bw�H7F�!�&��V��I��{Ju�Ɩd�q��@�e���K$�M����H��%�83Z1�A3�)t�ۘA�������a �;8]�r�m���Ui�7�Yz��b%�����	z8�h�gG��d[����G���Lwa,k�Q���Q��\j�����6��u8�S��zۯP7c��pdX��5�Iu�C;��q�b�c@������ܴ�Q��� u,�sy�&�3�G��
w(tg�CC�î$(`H�3��g��cj	��q]6u�IMk������!G�P�;B����%����u��Lbeӣ����q-�BI�!̣��.��0�-%��f�ȟ~�ԤI�sC�>G� <�^ߐ�v�j�>[(3�8)~_>}�mW6��d�<��;|ʨn��ˍ��O��j�������$qC4�˵�H��� Ez�����m$��c��ȗ<�v�#Ɣ^�3
�&�w+���|yˏ�'/%����B�`�频
��d>�Wg�m�A���� �*_S?�[�ܴ�_?<	vR�w�q�ŋ�����Vl{�,�Sw�[��I��_W�J|�_ʽ'�xt�W:�Y_�k:�$�O� ��褀�	n�J�p�e�$�E8��-��FME0�Eb��r��c����;`��G���3Yn���[����^|܄'S�-j��l
'�t�l���Y�n��*���%��)y�R�1ĦI~[�T�H���.���P��׆D����!-Ak��'�qP��G���������+���C�@�tb��;���_+Nk+�hal )�ئ�����*D2v؁����k���c>������P��X�Z��/�r=�j�zC��!G���Y�z��'�;¦:P��3����%�?�}$�v�ql�a��]�&!i�b����[�h�}�o�'|*mY�dL����Dy2T�\���WǦ���ޜ�h���td�8;l���m�}0�/�}��0�^�'�
��2�ؗ:��d�]�xo*�z�<$���0J��X�"kƯ�s�8^��b�W��鹞��I?7B�=�wy�{q����%���v�������1���p�@��Gl'kV��圞���[w��='�x��RH��
�\�4����?���((u�y�\t��^慲C�&�qش�Nd�� ��461|߂'Xg	
�r�I����d��`%��Xz-�N�WO���1�f��� �i&K�Tkny|�ߤ��rm�Td��+' ��Uf�ܔ�m�D�"��*��aH��5'uyX�V��J�]�AbJ�=���0������hL� >�<�[a�uG	�h��dL,P}��<\C���?=V��(�ӣ�	X�2Vaa�|Ա�`�|p�W������o��I6�V����G6j������P7���]�Ն��i��5�/[1�?�k�5@@-�_�aZ����Q����d�=Tq1&����Ш�%���[���XZ͇��KE+�Lp��[��D,l��¹�L�i���BK�m0�ϋZ��2����3V���[���xɏ�.bF������[�{{�X8׌)Mx��n�jw/E����uT���,9��8���_)'4=�g�)�G���cz���H�
A���q~8Ĺ�%\Ob
����qV|��R�|Hت����rA�A�<�B��.�+�wG���0�B�dt$EuJRL�/ƛ�?k�����J��i�Z�ս���������#rm�8JGbI�>��w@{(UkT�U�ӧ聟xi�|�v�E� z��ya.Gd�h\�D�+;}�}������h��9��LbrhUK@vla?�f�֣]�L�K��qcdOf�]�Z��@j�p���J���%��a�"�+&O{�k�+�,�V�|�x�!�G,ѩ3�\H�Q-*����X�(qٶ�ZK�cR����[�/p��L��G��|�~��Rf������v�w���(��	
�#4�ܾ��C��<N�"GΤW����{R:�^�O+�s���q��P灮�$Y�.� !�_�h�S���4k;@���6J�~q��h�����RU��S�]�w����=��C+�QsP�;��T�]�'F�*�h�7�/���6�D��xL�Ԁ��YL=G��}pQ��sN�^:w��/C�i"�.�E�u�X����35���ɤ�M���K-�b�����:!��l~���d"ɈGza�1���Pb4Au��d$�nh��q�� XHB��x�C��/�?(����ă�O�f���S����Y���	aD����5q{	��GNw����<��{L��g�IH��v5q�o�g���|3��*���8���"H��<-s͗�b�<�i�O��u�r9�ˢ\Zt�>�E��>䏀��� ����}bz}كG�p�����Eq"�#���]���3Ͱ�*�͋��)�S��1��B�E��C]�A"B��1s{����FdV��C�?P3�X`�#̖��ܩ~��s3b���������z��>^�1�~c/�	��~#��v���OO��wP����xC�q�T'GG~R�9��M�w�������Q ~[��|��L	�����7��A8�؞`w�)����G�����{j:�PKZ�&zلq�X���z
.q^�5x~x�jF���[�%��	�j���]O\Hc�[�j`@�J~�9'���㶳ӔN�)ֱ^G����S�"X����S��@�+i�.W�����Ж��A���>�͝�}ܱ�����Nni�.у�%�A�R�;v����B����Ҷ��/�-l�f���4u}2?W�hG{�薮�-H����
�O�� 3���nTr� ��������O�$'UI��}�ON��&>�aw2�	H��h1
f�X�*��f#��8�Jq�E_�����q������Z�5ԖvC&RL�+<֣�}�ǷH�k�!)ɂR���>�6."�g��`�~��AP9!O3Bx��咾b<��
rϓ��`*�9[��j<�M!�-���W�S�4� Eg��7Q�X�%�h�/�>���o
?�^{�wݢ+�%R�ۂ�D>�J�-�-�v�O;�.�j8 ձKi�2<����o�����p^:"��	�%�2�ܐ�%JAS�(�j�U�"/��'����r.(��<ܮK�ȮM��4�w:\Dv��������܏�翴G�f$�2E��AĂ+P��,A%�z�x��]�i��fi;�w�97ı��}�V���R�����0��s�7��I��f\�
!<<��y�ZJ*lº�ڸ����	u��b�r$�6}������&��¤B�ż��S)�z�!��V�637�[�`���w�_��̰���ڑH����*�r�uX�Q�6��̍�ҿ������I��y*}�:$j\^��\��%���`k:��6�꧔�$6o��;�&2@t�����W�a��ħr��Q>��{]�M/������PH5ƿ �zש���^5�u���A0e��
���$4؈�:/�J��/Yf^�o�#�t�1�cB�#8�̌�e��o�jf��1�[W���]@�E�cل0N�&6��x]�\Uߕ\��;�M��[c�	s���t��\_���[:%F�<Ez�vh�c�^@ ��$����n�FSA]qhw)��Mx����g��s6�5	 ��i�^C�&�����)��C����띉B��FY�'Z$�/9>��_)\	G�YF�A���L�2L����
Ux�Y?T��@�˱!w��	0���-���cs���0���le��Ձ�s������"K���e�����]��ZLw�Q>y�Ƽ������a���U�P����  p�B6Z������H9_��ZP��hث�?�WK꽆����6�QA��Dᓇ����W��K�W~�aw�ކi�������Ҷ��݅�ӻ�(,5L�~>4Q�	�*�̐��m.���%������MbՋ�}��H�OM�X}:�D�� ޭ� JSH�F�!������?g���m�9��Бl
��$\��j1SJ���6Dm-G�F�NϞ����;1�0�fw����N��S�w���8�*C0NLE�П~Di��"N�I����6Ω�f�����:��͢x�����<��+�T��;�S@b�%��` ��@I��DfI�֫��X�&%����C�f�jS��?�,�� ��̢	iD��,u�v��b�R\��Բ��\z�\=j��4]-��x�o%�QU���{gV�k5Ъ��QD����xh%����
�Ru<�k�������CwX<��qfX�����t�nH�sŀ���1)����7�J^���yuJ�se��׿rg��ڞ80y[/��&}D���xǶ��jh \㓠�Q4'4�����9ә�#����� Q�6�
aC�hCecBn�Of8��+*(~ԩH1'�-�T�f����-�#@TmM���%N;t4�neN$&�4��8J� ���T���`�6ug�S!�w�����7%W���+��� �調������5+������M�Y���qY��\������D�6]�se��o��6�����	k�*H��(&�Q� �R�8V�4\h�:!�u��Nθ�?�l�r\az)�{����n���ݻ,�'��_6