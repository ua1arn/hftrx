��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�����P��N�$n��̺ U�ˍc�� ��b.S���Q0a����
���`\�A{�Y;{�oaR&�-g5뗨"b�3z��ћ=E������896n��̹���)���UV����V���ɻ�eC�0eu@�wlG��`x�1�LR��1l%~��\�Ю�#�,\�xgl�'_!a�v�:����R���H5ڶ�I}�b}B/����@�*I)h�wϋI�*�����p���E�'�$=����G��z�U��c��}#��!�2=j�ܛÕ��N.�-������[x�vԵ�PK�(��2O�
����8ӕ,d�u����t�+�s�"��&�}�ԝ�(~���?�ŝ�j�����S�����r�>�\hW�Yv���ɸ��|5�Q}/]\Af���{?�mJD���r}΂�O]�v��I�r�g�����2/���6��n�i	��Kmm��~ĵ&�)�sܽ͐�YS�q��IȀ[��!K����C����~�����_��w��Q�z�}��W�<{�I}Z5(-��g� �Y���iW��S871o��@<��g�������g��%�Τ���w�|���!�X�	�}a�H�/��R-Pe?J�$	B5.��~JhD�(Sm!y�Y�1{Bu0��0�\j�����U4��������c�O	�)�t�T�+�Wk�dT���r���k`�dH��-�X�!:i���� ��*)ǛP=���ҥ�g����33��V�r���`�2&U��Z=�ZAƌ��#Mn���p�������|c��}Zv�� ��XD)�vN�w��_�._��7�$�Jt`�~������x�2
��=���j�t|�y~tg��r$t�kE��.�P���a`Kv��n���G�9RQ�����(^�ti��s/n���S�-�Z�W>��K��mIɠ��V�ҡ	,��a8��)��gM|rC���*u�c���-A�X,v��QJbް���%į|��lzw����S��A�����g>9��w�9�����(�!KN#Q �
~��A����Z7����RU��dң�"uޔ�+ �?r�P4 ���J���|*
��L�v����h���-0㮚	�' =#�NP��A�S�_lb��U��c�6���0�Q@�Q���(_�� \�����X�X�U��\l�4,�b�������9��]h�~��M&�q�l��rIHO�-�kD`�* �<��_|�����|�@v5x���q��8��W+��5W[8T0��l&	�;�=>I�#
v�4�>}i�a������1ͣ=��I	"�"~��Z����x�����F�F/ĺ�R=հ�����D�G�f
�l�k�!2'�tƊѲ�E@���¯wS�N�+�����, �����4D�mBV�c E����.qU��v�����.�BHFVhB�" Svi|�ȹi�D^Q��a1_�cY�@����rPwYԡ	�^J*B�-�6��g�]������1�3ד����t����%�=��`m���<�$�blK}+d�~w��a�\;0NP�v3a<�@��ţO�ˋ��㋤����$ԯ(��E �F�b�^ꨛPHk��`��_�+$�]�S�å�AEI�0`	rx�vP��4,����-�k��$�G��0�i "���^[7s�������?ᄊ�z�m�4׀@ea�x�_Ͷ�>kf�n#&���e��T��+%F#ӣ����$�.��g��~(	�2*�-*�M]Q�/M|L҉JY�7�X�d��F�\�	��͠�S��1T;4:t�ԍVZ�P��`[5����z:�}��j��x�FXK�g�>T���� |�����;\��8���>O(�sC��?��@IYۘN�3�<�8#�\�t4��{w�m)YN�C?���9P"E��K�u�#�-�\"��x��=?_4Lע0#�7�Ey���$
��r	��㳨���,[������@Rt�����l�pVs�g��2TʱsLNmM(Lgge����G٤hڧ+��O"�s$Ӊ��[e��%G�V�7��(b�M�7�����Ȃ�c7��֬�x�w������w�����7�v8�6d�/�я�I�T�X��Ò����l�� ���Xص�#�u���2}ٹ ɔ6�C����8��`�-���A�ldT��P��`HKG���]��%���7���⪻�̳T�ѫ�p"�өH�Y-y�'�M1�8��5��;'�;�-)�JwЅg6�ћ���]���$� w{��$%�`�4A�9�>x��.�i`z-�yU���ܗ+��|%X���2�gqfyG��`p�/�S���E� ��t�{��R��ee���'��-;>��`hr�|����4��X�h�a�:��"6��	#�����K'@����]��Ǫ6�o��ҧ�.C�J@/"�z2��9���\&ɜ��b�}��N���1���~����N8��+�!>T�n��v�Sݖ����ܪ���.z���-�6${����8Jզ�d�&Wl�>�W�S<������D��tC�s�a��qNd��˖>��TB��`q�V�O�;n�43U���NUf
�U�y��XN)���i���$�+_�i#^[A],9���b���m�Jp�*.��LC��^�Xdwu)�V'hA�TDK'7_��U^�u7�:';�I����U)ǡ��z�dw�(��E�9�K�"$̗���M���V��׍Ԥ7q˙�e���W7ӣ�{��H�\wC��1=���Q�j���m������[�pЙ곂)��p�9�H��&Z�z�j*�sW��]H^��\y
���;I�2�r����$�9���m� �F�+j���I&(C�([\����H�Q���"q��LX�+�j̑ۅ(�<�0[v���f�hM"�i'��A��q����T�W��i�.[���NpĊv��-�%<�ڀ&��,�`;����mC����Ǵ	7�ZV�X��[�-Px���++A�:?>
 S��T�R�=`h�ax)SR�W�=�T{�y�5��J��"�6�٠���iw��|̳v��J>8�c,`��bh����l0�zp�����Qw�(�e�����=(�z��-P���0���Bo`.�6KƗM-�O*o=�!��6������1{%�{/3�*q�}��z\�i�qhp7�p�?Uv�"���q,�P�W�����Ae* 8��!��˷��	���G��ir���փ��$�~O3fU�0�X�*���O�ݿ�q���RE[O����ܝ����1�WT�������k~W���B�Tc�C s�b+����/~�w��r"8�����hG�����k6H!�i�{�D��ݛITN��p!�,OM��4��H��1VŢ�4r�:�����Մ&�~i@�~��>2��E:��tv�S+8]�^fӇ��a��z���[�����U@���qG�˅���.%Ƨ<�i��mU%�	5��0��v��<I��Y~�%x���(�2����~8WZpa�F�U���� ��I�N]�3J��x���Gg)��w�ᨖ��ѻ/6�a%Z#e��k���%ea�>P����ݱd��$��+sՀ��d�<�v���x��@Ѵ'Y�(��bV6
�D�m�'W�}�$
��5 ˴p�{�J?MK���^ 	�[C�ʐJ�>ޡR�R<�Ijl	�b�.�L=	E�~�[��QJY�N	_�Ta�?�?q��Y_x,���eD�����O֫I��G)?cu��X}/�)���.A��+�u36UmԹ\;Dc��ﭳ����
����Bh�8;_ ]��B����{?#�5���$���CI�S|���W�J���Q���P�|.f˱.x?�ي��"�{j!���&$<-ݔ�Ir��,�X�*bĸ��a�CXf��l�I���o��NI�2}d��|p�Wxz�:[�K��o�Q�G�^):Zx��k�u������a)y/�jX��Dm��%$z�����!ry7�c�Niy��[��PK�d��J��%!�^��4U����S0��Jz$A�� n������@�̗�Q&���t�kM�'�r]ur� f��.K�/���(�F��	Av��t��(��CJ�b<bY	m�$	=FC������hrm'�Y���̼�X���$�D5��������rg��1RPˢ0#���D[2������xέ�<��0���c��4rm�H����r����n+t������ۢ:K����﫛_{dA�į}�$	�~H��V�3�c!�-�<�_a08K:�&�x&��݌n���F7���I�S���4U�g�\!�磆���X�Q���nT*��(3����!�H
��:}F��q�(ﰐV��.�S�ёe���C/�h���AQ��3R��lL;)�^'��+��$H��?�9� Y�γ�"(h�{Cz[���}Z��ֿ��/��C���u��{�)�R���i�/�{�z�E�_{�g��U��!3����b��-f�����ec�����S�[�>�/�b���&��ɥ�Ϊ�-f�� �NW.���Ӣ6{�D|���\\����|����������L�	I����sU�{<s��:��u�}�z��{�w��m��&���M�[�����?����d|����H)��6Cǅ����W���9�K�4��N.RL��W���ji1��2�۴Oz����ţq�P-��U0yV۫�:d����K¼�� Nq�к�xc��ap�փO�^������O�֝����5�X���.)��n�%B��<N0�F��w��X��'�_ؖY�9R����)-EyRXUD4�B�r->�<>U��2b�����O{І$zIu;�1l���\��Q��zo���B��S݌,����X6�g�v���+�� �tk^����Ay��:�{Gj�<���o����mZ^���sg�O9CBPƘ5��ԫK9��SK��æ:��j<��XPS�<q�{ò�/R|��� V�g
���FJÂf�²cY1�6�'(�.F���Y���<�k�fN���$v<��.������`��g�L�3��X<�Wĩx�}��m��ϸ���#	����}�O O{i8�[&q]��7sE~�{��4�@y����k���>��J�=���jG,Xv���O�OǞ]���6���w��Bh%zO!�]��]p2�y��
�'��s�)	�5Z]�`iq┃���"tvnK P�nݩf�Ǒz��b�W=gX��fc�F�%�����R����Sy�����F�U�q+�w��h�8�-�֓v�8���pm0��i���r��2K���fE��,W�����ƪ�Ko�HPw�{�Ts�3%���.���0���óI'(B���&����-HQ�@<B�H^V�K�
{������Wu+΃��$Jv���Z;2Ung�~y��;���Y�p���ue�n�&��]��d�Iv�@�VBu|+8��������h�R��y����oJ�7hM��ws8�`^��د�Iw������*T��B�C�t���U��M˚��� �jKG&�0Z�=��󗇈}Q�&�Bq�͈����"�vR+0:��鷉d��n��R����Pڋ慢�������V�]P����Z���4�}���,u]� %�R��T��k?�-�#Q3�p�Z޹�z�7l��aų.�^�0Ě���B���EC�w)��-ۚZYGȆ��@O���W���y��DS6�)ra�!��}��ta�JQ&r6~��DN#�Dq��/�_i��2w�)r4	LG�I�y�:c�ڇ������*���{�g�R'����q-,}n`w�ڳ��Ko��Dʿ���b���{g�β |i�5�ӝ�k*_���7Z�� 'T�h�﭅`7���r����u ���t�#��ݩ��)��N�/��y��MĂ�0�A�h�Sc��|~I��O�h���L`]�kx�bȚ̮���!<]�Vw	�<��[?a �8��-�D��"C����Ҭ"Эd�7x��J���\,*dOe��Za�y���HC��m�/��b�l��6>�a~�\�#��'��(���n9���;��=�G��:����ě���k7�xmα�����Z�o1�`�gUI���ћ폐����3���?pO��5j��<��JO��⅊� D��� ̠�洽�z��~�x�	��n�.ϩ�!��i;��q'�������6�}��� 7��qARW]�r�8a2>E(=�����������N��\��5�ef��s�����k$yf�C�LvDS�)"���f ��O��fkK�����>|Ú�}�4I*1�D�Y���Y=��2}g�>�͓�T,����,-GX���s��f��=j�eI{絩���YXx�