��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�S�T�;Ϗk[�^��_�5�
�V���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:��׶��{�*Z���H��ea�8���*���g S;'N[��I�]P*m����)O��Ξ4�"�\�� ���K�O�{��׮���^�ן��A�ߙc\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�(����5�2���[@%����nEA�V���E<v��9�ĒTC��0���۞�^�� ����C��H$�ƵoB;sѱE�ouJ��p����B1�o3(�'�"̂����b4MI�-`7�(Y��;(��Цy���t��k�8���҆�|n�����|Hj`;U;�c=���)M�BJ�Й�m��/K5r��!����%�J l���&��RL�a)r��fI�����,�%��a����2��>҅eB���u���;��I�6r���ScB��\�~�q� \���T��U	�1�_u���V����*�^�~ì3"� �vm�!=�y����h�}��<]~8+|���g�S���!�<o?�M��;]l��j�z�	��A�b/���"��y�s����o�k�8���҆�|n����e��m*�~^T�ɴ�#���3J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|A�־���1�9���1� c��(�U����	x]̍��;����8�t`��g؇�"3��
f��:�%�+M��m}on���b='��\�4�s��{��]Q���/P�Q�=�VV}��ԏ ��	Y�'7�~�MUs �Tx�B��ǩ
����z��ee�:�$�i��Ahh](
��x%i")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�<u�<�.�Z3��a� ��l5��e^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEA�����G3�7DY��SE���ƪϤ�Yk"1/���%	v3־���1&����k�+}$#�s�'b�t	�U�lZ�K��>п�p=	�˳͠m�xW��"7D{��\�v���4�u>�[�9q��q���U���g�,P�nZ鎬�����,���
e?V�6IWJE�r���秹��ч����=ў@'���Xw���RY�刨Ψ��F$��O�&��;�L���9�D_�3���U_�+XٹC�ߠh�N��B�)YN>�4�
��o�M����a�si՝�3��Q�B�1Y�ΊS&}Z�F�>"�ѐw���5�W�u,�%UU��2��{i�X�x $}��}�<�W�C%�*�JvW(�%��b����xVg�uP.},d�z�m�~��Z�H�(�*�b�βł1Y�ΊS&��$шe1Y�ΊS&������'l���u��-���E�0w�m/����;n����開ϡ!�����΅��u�Hu�@}H�X�6䯟I;Fk"�i��\�v�JE|Q�R�hbvk~�#x֥�Jamo�/woP}[�.ᬵy��@ӌ$�Ê�8!��vp�P}��O��>��Ӫ8߼
�d4I�<'}-����_+b���z�d�X�VM�����a�"e͉�Xk_�0��'nU	b:Nn�|�",ӓ64�)��8z��uP�T�UX��v�^ܯ�~����pؖ-�/�+T���u�I��'�4��,ޫ�^o��>n��rs�i���\��_���W�A#�q���U�T���u�I��'�4��,ޫ�^���D����q7�F ��W�A#�q���U�}�LYO���s�����1�:�Ω�S�T�;Ϗk[�^��_���+R 
����L�]�b�֘m��+��$|��;D���J7"�dÂ��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��ly�(&�N�����B���0o����T/{$m)mW�/��)�-��DǷe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I�+�c��Uwz�@ʶ��辐�!JHn��z��C��ྐܼ�\�v�9�#=�8%�b9���J���z�my±�sR�{F  M��va�{����PD}#��ůN}�m��{B���T�D��\�v��8&���I���8|�L�*�g�;�k	�oG�� h�ҩΣ��n����-�����y��j��k\y[P޽��5 cd��#�xy}�����H4 3g�Y�T�:5A��p��jVѭ@�y��j��k\y[P޽��5 cd��#�xy}�����H4���b�%3�;b�-�2��;�P�t�5��w�w:�;�jmT�#q�P�:땗� h�ҩ�p��xs�S�*
�DWo$ۯ}z�| �8b�9A�i���Y-]�\^M�Ɣ�	��x��ݚ�Н�
ҭ�3���#���1��t�Q�n�!�&}Ji��6���l]�a��}Dq�f��5ߧE4��HN��R��bP�63Z�t�y�"�V��5M��z�o�*� '�!�J����ϩ�Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����m2����H�� ӫ/��m�Wq�
Z*�)�J[x�*��rC3�8�c㚂�IB�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a%��b����xVg�uP.},d�z�m�~�.4g$�co�XB�&�=�b9����N��a'��@��(5-ˤ���k�˒�����j�'l���u��-���E�0w�m��<�mlo�2N��n�=U���iAe��Y��)�?Z����JHn��z��x�f7﹏,���D��a�si՝ӣg{��aDeq��ҝ�r<�n"��g�LX�,T ��b�FP&���rS�h!�`�(i3�@��O���Қp%�0�ΩyO^~��M����A�m�(��ڽQ����2N��n��t�J�Yy,P�aw=��E����F�_����ֱ�q��w�G�ïWA],S����|:��ͼ�\�v��8&���I���8|�L�*�g�;�k	�oG�� h�ҩ���D�Ώ�ƅP�!�Sbb�����@|����r�����L�����U�ჴs3���l�c�5ߧE4��$�[��= -|�GP���*y}e��p��G]@w���a��G~�= cZ�-ڷH�%����@|����r����~Ps�Й���a+Q�� ��s�gJM!�1�� HN��R��F F�E̠�i7N�_�z*K��I4��欱���j���]���.��|#HK���v����`!�;��!A2�WA],S��o1s)�u��r��o|���P��3��/���WA],S������=�՝� s�#���k$ �<�I��y�fe����~éޝE��Qfĉ>99��A0ok����DFTޱ}b�g3�UX��xϚӬ�5n��/0�E�i�m}640�RS���$
�)N܉}�B>i�a�	KX\�B� �b��֭�h��O�Q��ǺΕ�A�m�(�O�Ŝr{= { _Ta�F��l���)�4�����Ὡz�*<�����s~��!��jVѭ@o|���P��f�Nd+l�Yҽ֗��Ǒ�o���D�Ώ��V�:�R�;�P�t�5�37y�����:����@��%/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!�_S�t�Aju���lWg����ha�`�2G]�Mq�}��,+$\�M���5E�[�c}�sX�>P�2-i_�	,JZ�!�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�NilM"�����iM0�3m�:3��Տ�L� $�3"���N�T<1(�d���Mo�~$5��_������"~6���aq�����4�k�߻P`���;���N���M��A���va�{����2����%��/q|��h�ӵeoQm�`aĉRW�F��F�zL͊�q���Z����p��J(1�:�>�̸��oJ(�c�-1F�]�q:��c^�Զ]܆�����ң;�f����~����y�Zk��~��6n�L�%��/q|��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xB).V44�o�.ᬵy��ՙ�3Ќ�L:(�
�*S|ò���
��_�����k�79�����\�v�%�M�5&l����I{6���>�3���/��¬3T���&|���BY��l��=5;���ip>��<ug	h<��Q�R{�lp�q04?VS�����ud��%BJ�g
�zP�w:Ec�[�p(	��Q�^�y�zL͊�q��j.��?�Uʚ7�ܩ�.fOe	�o1�ֵ@�3���/��;L�=Q ��b�FP&����҅JHn��z��`�+]���e���im��mų��n��Uʚ7�ܩ�.fOe	�Ƞ�d�P_�n�To�[�}�~��l�}`V�u�6������1�R+-h]��.�{+�&f��w�'�4uB���u�~����J*�Rs�0K=X���d��J>�߯�"5�o٥����Y�JM�b��v݋N�����7u7҃Q*�6������1�R+-h]�83NI�����w/,g{Y#0����l��=5; �e�B�R���>_�4uB���u�~����J*�Rs�0K=X���d���fx'v�ao.\C�k��|��-�Vc�$J�{�����~�=��K�I0���ԏ�.fOe	����4�l�>z�Vg.N������[� �I�������m��b��v݋N��������џH�5ߧE4��?"�����2$%-����y�����=u~Ei�"2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE�7�0}7��k+�=Qj#`�,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�Ia�6~n!5�$��fP����E"�T��b9���M��A���D]�$���k�1 �O�o/��T�n*�N}�m��{B���T�D��Ψ��F$��O�&���e�JP2Ud̞��>�1���t�<���8-|�DOYZ8�%QQ�{��x/��Qu���%<i�LE� R1Xi��&\})����K����J���y��j��kj�����N�_9�R�5;�Щ�j#/M��\�jX��u��A�0�Ή*��a��Ɇ%5�����{��ü��O��b��֔N���c.�'}-�����@E��=�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��0���V��C�qҢ�����N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開�Њהt�ȳh�L>sP"G�wk��a�S.l"�S�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3���/��kOT�i7N�_	�z�w.{��w�_��(�6k�4d�{j����·/ҳ�ϾQY�u��A�0���򴶽!�y�"�V��5M��z�o�>��U^[U�7�tW-�J4p'�>��\��:��Z鎬�������(���w�?�b�>��]�!��=���W�N}�m��{B���T�D�]�!��`��j(&�L�i��ko�$ƍ2���lĦR'cf����T�x��QU���^4��y��j��kL1���oB�T���I�!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW];��e�8<�V�Zs˿�}w��ea�8���*���g S;'N[��I�t��ݛ�