��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^�}����}�n(n��z��ncf��pf��Oy�˜� W��qI�ux2�LdV�ٽ�X*WC�D�(f6#YX��V�]�u��:�	
��m���42�]�&�e%#^׫��M8rt��@,,��:}��Д�홊
�7Ec�]���J84Qn'��H,�$� �K0m�ޝ����y�,�
c	U-R�kL]-�T�
�ϗ�D��3跣H&�?�5��ƾ���3���7_(��i&&��<���K���.�!���5,P�IVWh��:C�/�W���ˑ܁/�p�ّ]�#��M��όu�2'��W�wӾ�_�z�,X����܉����R�q�3� �ɫ�3I��ND����������8�{on�:"|��*��'N��b �z$����x4���it�e+��H�%|կ�u�66�Y�klX�r�z>��#�GA�"���5�7�(�~\t�X�[P��#�=�վ
�id�p�[�R������׊�<��<��ľ���k�j�L�
�l5�t|D.�K��]��[O�d��~�ѷ�FN4@�V�h��>�OD�gt~p�Ӽ�R`��մ'\c"$��?!r%sB� �������#n����� �pҍ hp���ʳ`Kl�������Ŋ��<>F�p���;I��������F��[�#�@��8���ώ �*,�&7(�z"�x�.���9�tq����b����N��p\��+,raN�
� ��d������lTp�e|��5u}����пGe�<��=YҒ��}i�bPH�;���ט�-��e�#�m��N>�n�\�ݟ�ͨ��IzLkU�U�����?bzW�����g��3���D����݁&i�nF4��%�~�eҶ2�K*���5��`�㑅��8���
r��/l��9�LL�N� r�=��Ŏ�;&ׅ����?�m���E@��������6����7������|q�JB��Q�vqŴ3f'�J��rB�z�+e�r���7��2�))�Le|�|����(6`�l�0�L�{�0��r �O�8���(�t��ڗh�C�
3�%$�4&��Im��B�i���	�)rl�-Q���U̫����j�[p�Ƣ4k��E!�X�OOIZ�U"9�l�^1�$Ю`'$L"5Q���8Dz�'3!��t���A&�K�]����Ekf��q��|(�s�ʣi��Dw�+��85��8rz�ou���D;�r_I�����.8@�GY{���u��Ġݧل�I������jZ,��&@��������~��>>l|:9
�!��� �gFpm�^nm`U��ڧ���~��~�Z�����'t���?�����ñX*�8����rM�f�ˆ�4�I$Ӹ�%�K�N�l�,^?h���ڄ��>��F���Η���*R2��̏g�%�vK����&jO�G��N2<d7}�[v:�漅'�^5�O!�Bb|�������%m=�]�J^6'yq���g�}=�q��+3-�Ef����F���N���4j�B-<"������fڻd�B4#fY��:f�
:3�t��S/7��G�V9�w��+v�'��I�L�$î��?k�B9-�X�Md�VXF$�Pʄ9G=h�F�wJ���\�A�5�$��.�����#7�� B��k�E�V�6��V����{h�J�9�z��w�3K��
�Oc�8r�0��y��Q�~T���i��ދ
g>�Kzڎl$�:Gp�m�Å���׸�׋��i���v6Qk��f�E7[�<P���&�pG~ԃM�.��JV���6"�5��y@.�Ho� �HsX�j�h�{�"�iJ�yq�X�.ϱ���o�f��&`�[�pΣ�hjEH�*_cK�[�NX4L�� GMi�R"�� ���Or��@�\���+6v��fWk�����n�`.�U���z���8�1?�!������LU�o�(t��i�_�SG�G����ظ����D+�[;�A
�
�^��g3��֬��BH�uи�H�]]� R���f������ܯ%��i7����+&c�E�h�m��}zY��A��l����,�L�O�.�p�$�-����`���Ge�5#/����־	���4�;O#�YV"���0����(��.� �X�
���v��"�q��/p�9$���+&�n.�oǩ1?�Aa%�065�()��hI{t����T������&d���O,��.�lI6n��.�4>72j&���D�����o�AJjf9ԩ-�׿%��A�f�]��nE�k�CQM2������m'��7�K�I,���ٔ�H�9���/Ε�ݟ��+�����Ώ
_��b�6��8/�y�x{i��t4��v���E�m�����gy�e ���U+�^xy��O�F��MxI�ޖ� kЊ��r������Ȍ~K��x|�ŋ`V� }���>�Q{8U/��CԾ�X�����U�)���bT� �@���t���yt�'�d�Hk��Ш��� j���O�Id��6o��jɡ��Y�渠���A���iO6�#2�����B�ʪM���D*��ße�N����� �O�2,�e8؅����Ө\j��h���9�7��gfn.E�+�)F1�]�q�X`7�Pl�t��B�����8���3�`�^5[��Wy �ɦv�Ώ��b���"��~�[t��t�=%���,k�W�VȜ�)��<H)��u� K .�sh��S��j���-dO�����A�n���P3)G��� �;�m0~��%���t'� P�3�OA�m�b�j6���$á�BR���L�L���O�mz���l弄7��C��dIi��]	��@tѿ8ɻ�{Q>s+Q�z �����;= j朲,��ȳ���G��:�0�C����G}�QĊ�UF7��|8]�\^�6����g�K�ٚ���T̏�Z/b�ypZ934e��&7��.9i6L��c8�N�vOׁRP��y ���a����&{�.��Q���R4�@8�tH�E#�kH9�:�r�x{�����E%,xm�K��/�	Q�/ͷKo��8LFZ� ψ�%�[�?� ��������/��rk��d˯=�z�X�_����Jvm�|u���iD�V>�􏷯-��S���
s�I���H��������1�a>ϱ���Rǩe��� �PA���Z�"F_nmc���V]���B�Y�{ĉ�ƹ�m��=EDպ<�p����Fm��z&y
%��b������7z�����C���U��u�.'%��}�l�W�ehlMf��|�[wZ�.aKʸ4w�������FV�n�����Rs�P|��jA5���O�&��e���Ӻ�G�&���kWPU�P64Q�1���ͳ���2�cf�2�҆Z���y8��i��ݛ^�k�pX���ǌ��)H��{�$"AGWRf�����35R��7�E���>_��t�W�/����6��L�I�?��p�9p�$���Y����5�V��5V���ȁDh?�k��V��1k���	�۱��iu�\�ن_:`��6G�擐z����{v:r�;�jS}�1�:�T8lPP$]��M��p��9����I��v�5^��<����D4_O����}M0��7�J�E Ng�N��Y�xy�7�G� �$�YT���}�c�mط	$���(ʻŵ<��1�$�'?Y2��B�T��~q�H�1K��H�!o�O.��&*��|1A�Y>t�]:��-"q��*��g��,'��O�F�����m�����א�m���
��|T%�f�>�h�K����5٫$ȍ���\g�"����G]���{	x1�n�g��;M�EI�/��<N�d�-)K=�6�+D���I���00/�3ڟB��ψ���η��+�yJ�hn���4l�	r����-2L?���Ij���2I׻�z���ѐ=c�����j����=cY�c}/ǭ��c��$�^Leg;2�?�C�;�~�����(�@?�ޟS�Ok!Dr��O���}���fUo�_��5|�� ��o>L`%��z�y0��/�2�$A_F(T+]Ch;��Ԯ8V{� ]�ꦫ�-f�\aرO�х=�����OI�'<~Gvj=��5�������3R��RK�`$@ݍF��s�BRJϗD�s��U�1�@��g���gdRZ�S�'��Aq���i��Q������M�%	ӊ�)j��n܈Ψ>��D��zH����J�XD�u,7Ε'���hFg��.�����ˀd���m�L�����ƍ� i{[U�j���dѫ�wT����u$��Š�[f����n�T\C���>?Wp~�i�(�*�����u�y�3�zt.
g:��
1�^#��ab�e���⬁&����8���N��5�����h�/�?z��N~�5��rX���y�{�	@3$|4��b���R��s�ޒ��A���Y�p��ե�(Bw�7�^ �p:F+<��-d�[
z^�9��@��yy!xo�J��Q��Q�=Ta����eQ���\�x�^�̣�caqo��Zߺ��(��r*� �c�ޓ�ij0��
u� ܙvȩ�W�;,�t|	N໇��%�K����~oyXA��FP�d�|�e,�LVY�ha��[n{"��
�`m��oz�n��Q\2���)�V�R*V��<�YS�ӨjZ��;��6dr߉�"-��'����*��^,}m�]�?;��A��<l�ci~N���+�X1����f=�4�utIJ�~��V��ogPA��Sq�3,�A��^�&�ċ�nf���1٭�w�m/��s�q�s�=(J��9�G
�K]>Y�4�&�TT��MLs��*
�4��z��-z(�R`�����S���6��'#?��$�^��ݩW��CH�J��=��>}D��=���?�$��7���18O5����w�\D�"[R�d�cEZ�Ll86�F��܌Q�Í��m�ce��M�D��g73�<֕�&����tQ��>��h�"H�Z��(�X����D�D����sm�R>oc�?w�I��H7CR�F��W��#�aN�"gt�T�o<[�8�AG������vS�C���T߬��k�4��1ƛ��IfR
�����*���edx�����眼�^� [�UR�o��[��w�H�؋��\���d&��1�b�e��.�C%���� �XOm��<H�M����fo��~��3��2�=�\� :���I��巈[��J<r��&U�e|y[ ��Y���A�豬"?����r(�U�Gyl��]�� s�u
kS�� ����Ckp�SM�ãr��pe�~gN@5ќ1w�U�UrT�QAF=�	�����;h9
=e��T�&��ZR�����^B�H?~5r, ���i�4���\/ʽ�(JfH��*�Ҕ�sK:�@�3Ep��]_Oso���7��ŋ��xy-��gp;��3��R�]dU)K�b���SَeΫNI�R����3D����%FҌu�)����:��Pz��В3�4�{�VM�8@�Y̥Q�ў��=H!(�N�f���xO���?b�l�j�#r�A�Dv�ES��B��t;�ҝ��oH���_�'X������!⓭i�A{~��m�ڄ�a����͎�. Ъ""F�����	��?�$0�$?X�H�I�21�/	�o`��r��`�(�qr
��!�W'ϝ���%+�I�7;��k[������5ߒX�P���87�@���l�:+���jC�ʕ���o
<�  �ʵ���Z�� ���r��uf?Vc�ɜ�7+"�74��A���5l�G�����Y=�$fwb�2lR�.�[y���'���7�_��'ِq��7V��f��c#���H���oԫ���(���C�`��$f���5V�t�$6N�D�M\�ω2������ɱ���Zķ�u�ڞI�?P�	S��3�Y���+n��Y��}[�+�C�k����U#���ܯ|n�P�Qf���~�]ЋI%+W�Ar��ȣ��t���p�)��,�y���hl]��&��BS
�n6�s�I�m�y�˭J=p��>�]�\�5J���h3����rH�4�󥘜h�_��~t��fE�@�<0ɹ�5�a�x�6�LhEʞ��d:�~�-I
��o��XVۥ�ʃ�yb=�d�Mr�?�ǿB-Qj�nZ�q�Fv�>������}�״�e8��/C����_��������W������F#���l��3��_��9�l�$z�!^6�8��ȫ��I��\��H�,4�$�ؿ�X�/�\.T,?y�o�O����2�.���A8Od�Mjr��_���!�-�9���%�^����zh$l���p]7Ŭa�	���}�<�y��<w�����50o��>�-���̘��2�/>IrdˀE���;�~���2��zx��n��M�iA3n'0���|���,�����7�T.��D�����D�z�;ھ�����N��n�d0�p)7�(���4/z<��|k�:��l��͂�=�n/#	�����3x�ãv-��P"�Q�zz�J޿O0vΈ�[&�G��t�zx%�B��A�U3Y����Z����H�܅�Ia̡��ڶ��]�H�ӍWe�t9��p�=����z�n���n�Cz1̻���zwA��Ex����p�+V:��������p���夝��r�|�;{\�]����U#�m���j0��NN��(��U$PPZ���o���0Pv�[�B��3m����Y�-�h��w ��/���\�����Y*)��c�D�Uy�a�@���m%0x�
c7J�4*���^Q���i�6����Q�T��ku��G59�ȟ(砫�����i�id$�_��<5���$g��F9i[ѐ�ohi��h��T�b��a�X�.���'[��AI��\ၗ'�mA
���y@r��=$���&vB�6����ꘕ�7���6NzI)}|�������_�O���/�=!W������0�SKk���ϼ>�:���C�����eu��}^�偄zd�ʘ�B\�?�A�K^�d�!�������T"�oaN�l����A�b^ݼ�
٨����/D3�d������QƲ�T�I�����%�@J@).�G �&�׎lq�钧u�{���:�����$�7X��j(���c��zמ�ĭw+*ց���
�0�p��S9,���~�:-:p����m��@��I�?�Q$}9~�������O��Ǝ�`Nu�h;��n .*�S]�S�V�p���*:O$/a$M�l�̼�<�H��y:�5�#|��Z��Q��g��sz�hӔk�1�?�5j�J~GU����P���c�h��g�3>��g� K��\�o��d4�Xt��tH���BBih*ݛ�!G�c3kIɔ@G�@��^Z�`~�0��-jQ�9c�+�� 8E^Ҽ8�����&�[r/NCxz�ѳ&p�2����⿯�s�Q�ν5*�H��~C,K����!���D�A6�K�E�x���)ݔ˂�J�� �H"�0�r���i����-/G��������K�J���q������u+d��R�dYd�3Ej	u�k��F��Uoj��|'3�k��9�,�	w<�!�����BN�7ޯx1]'�r�	HU���쩤�~�CP�c��/�b\�D*�enm�!֛�Xb4�������>�����:'�6�{�0p�#��<=(U�r��I>�o�Ɣ9)3����
t�Lە_�N�����ԒP��7�,�L`G-��حb��&���i������o��]Z��ܴ�_r__��K����v����>?�x�h��ΐ�r�7������6��I�7(ڐ����
_Q��G��keٗ?��8\�3C�BD ����3k�`xOͶbtzj��%���ݹ�G���'����o�:�M�s?״-��ޠ5[7�����Rc�D[:��!�R��!�KX �¼8�}��S�`��<��fؘW��;�L,Ɉ��%)�lia�K��ƧH�	�H:V�/���`ʦiq��>`�Wݛ������ƍ���2a	��=xM�^XB�K�P���I��u��l�+h�(!�ٯG�Y,��NP��M���mGLݐ˔���eqC�Z7����4,�ҏ�zB�?s�ϧ�E�jG"#9�I�O�8yK�zو7��eS�G�vi��fj�nî��Y�� �F�H�7�#Z~�/"l��ϡ=���O�[�	ժp�{1J��I�Ԏ߫�@z5i�|�M?a���!{QɅ��̍!�;{��h$z�Bc��(w�A��<P�
�G��#+�~���k'`��q��"�=u�<����=j�Ê�ZXM�	��L������/�������f4�_��.zu8����Xˊ�Yǧ}��C�؋CxK`>� ��@�{�BL�&�O������P�������C��2���'�)��>+��b�t�
_#k���*���dgΔ�
Y����y��:ʦ����ݼ�6��~uS-f_�ѰK���K��i��IS�J��	���f_��q���V�7�]�n��#�%���V�j�#'s���RΡ��i��|f�J�$��K&�T�r�T�͌\��kv7�@U�ثq���	{�T���V`h�s�N����K��)���'�탧��Ӓp�K�=�ϓ�X$A�ah��kk�»'�Sӧ�rM-N�"Q&��Qɋ��pM��?	�V�7m��}�$l^����WT˕~X�Vƣ�(��}�4�  | [eǮz�Q��q�����r_�h����[;eF�!či�U��ܝ�)3���I��&��i@\�s���-��C�����Pc�2O��H��w�p���S�p�pYQ��I�(⧤}���e���N
6��D��N)���[򷞒k[�0�$��gXMg ~p����t� �'���/$�R[���0?��c��cK����L�o)	�0B�6�Lk�E����k�pDp����:��n6��}ر�Q��C�OQ����Ӧ9�ͩ�N�d�ǵ���8C'���6��JNw'�	�U\/�~�'��G��G��;$��}��'�{�6.	����O�o�G*�g��iN�������5Y����F�.�v,��N�{fᰧOq�UkyQ�������*���y��'�2�����=as�
R+��wÑ���n[��/0��x-b��Ъ�p��k������8�iiJ��|�����V��԰
�s�~Q�bDg�����4ܔ���܈^��ZD*�	�3.�+��Ual)���J#Dv̰�L̫ߐ�X3��'�l���]��"�MU�p�<��G���1#��Sm8�IZ��;˓��x-!�9��)�
���q�MzY󧏃 r���j�cA�$�gҎ�x@��T�7PH���"|Uѣ���|�Є@�k���X�6���/���.��g1�r���a��}Ɉ�$��:P7�y�f^S4@IX*C�=d�r�Vሔ,�Z�S�I�H��"gL��ZQL�����/��0"���(���%�i{�@�����&���(���yiv]����3!/�Ȼ�Ѱ ���Yꇙ�-`��sv,~	�z�(ҳ���JN:���s ��oU&1�h�d;�(�9^(&u�1�r���t����c�7��~�C�ʯ?RjH�Ë��t qM[֤US��ں�iN�z�V�N��	�x]ۡ}:j�71F��m~)�}EGMC++PU�x�G��u�{7����]jƑ���$�DC2�=���.��گ���n�z�8�yv>��u��W]�Y��h��ɛґ�X�o�1hZ+�j�a�RB�]����膇�=��@�>�c�K��F����^�=� �����zk�O�N��Xk������N��&�)�h=�C���4�`־.6��{ل��TNqĦ�u�8�W��勄��m���I��=�!�)s�N���]����z\.2��.U�`�~��;�w�,��l�9�~	1���|Q�����x��-�;[A)�]l՚"+���S<t�G��γ$�[;8X�:�L�'��,��ŀ�z!�04�ZC��B]L���<q!�$�7g<�B̕����I�TMns�3�,+I�ظ��I�iG�|��{�BO72��w�Fj�Q�YU_��zlxCp]ɋLU-��L���f��ӱ�V���"�?���V�0-�#v�1�OqJ=�;�P ��\nC�>q¶���M���+�c�o)7�6z�a9����88.��h��YJ��y3!~+�}���PyUU�g4
n���5,-�������7H��L� >��J� �M���U���
iZ#3Iԣ�N�r�<�4�����1^6__�X���D-����=Fʣ�]�$e�����C����R�%
�����@�/��wkp@�u���!�2\��F��@u��:s�.I=��e4�b͛^��Ó�L�D�5ړ��# �ia��T&4��Tp)���wv�1�=�?��4K��iu�BORN(�3�2CHI?��#Bgu�?�6�K��U�)�WD=y\�c�B��'��M ،� ܗr�,���b�7�����B���m<:'pH�S;AOs4�#��%�"�g=�ٟ��9=<�8k0#j\��2��!U��5z<;N����e��:u\͝! f�V�1W�ɀ�WG^��c���KN	1ӊ�Б���-�r�(�n
OBvME�ߌ<�y�BeĦM;X�j���E[+��]RE�C݅��C�{d���I1�"Rc����VȪw��yG��`��s[�TSƳ:�uS�E�.��n��L ���� :D���.��Tx�搏d�w`:,<�{�h��7г��~k&N:?X̆���=q �p=��9D`#5Ģl��<����r.5�2�F3)Bj�3�����#�F�!�?�P�o]ג��i���7��z�~�3*���ą�%�Lujv�� ���I+�ʋ�������p?=W���ޫ
1���)��|�_h���i�Dy���fA��Ga��ҥ<�.��G; ��qa!��7�i�>��Z��!A^4aA2(�av�1bm+��|Ԟ�U�*)�DpΚ&�Gވ���E�ء8
�&�cʘBv�z�������1��r<Vs*0H�{#�H�L+6m�����pr�ǟ���}��WQ &7<-"^u��nD/�To�%hd7���j|�ʹ�Y�^����j���׎l9fKoqOP�Wk�i�d<d�;%��N�	(C�N6��,cx���b{��	@�55��勤����y�~s��
�*�J�{ϔyU╈	�f�&�6w�X��+�
������[Y|�4n���&'�<��֝��+������L��:�8_���xnȮl�ii_�����"L��+�?EvA��;�2!0�i�t�x�7 �g�|uW4mc��A�)n��S���tP���a�8w�����}Z��K���Ͷad�|�ڸyr�l�>I�ˀR�=�����R�j��)۽�����:�����y�����O}���aj	��l���o,
̠� �������Q�:�]H ��NGZ��!]�̑�L#4;���i�&W��@v���]����x�P�B���^��桊����8����Z��6����o��h�"�:o�ԟ@����',{�DbK�zD������A�F��\�ڶX�V��|����Vغo�@����E�}���ʆ�a�bs` �?���� ��g��3����t*���t(w��&裒����K���A��zjN�����TY�p��}3q��F��f��������P����Ko�Ǭ'������E�-���	h+��'�U
�4#��-���d�ԀF��5+�2����G��:�-b�74�8��c&*�d3���"~ɹ?k%�����Xt�A�pvVf�KT�Կ�*c&��+]ҕ��|�������P�ڌ�5�; �.P�~CJY�Ak$�j�@��A=�RM���]ke���ETW��@)�?X�
r!�#p�1ߔho�	���sE�lW_��&��}�d���~H����Vԍ>؅���d\/���eX�������W�t�hz�K��gL�\ퟤ���s�	����5y^���U�����#�R-�q�p��D��°���,�1�Q,��'�@Q�.����vI	��/uTs�f+d�{� 5�/$޲VGb���F�=1EG�����'B�>�T�wR��D�6�˲�~|�ݳ��#� ���ݖcVzu ��m�q���)����넆D�O~mǎ	(�E)XYw۾�7��)j^9�+�.*��`#Ho�c��K�m�m�)H��q�� ��{�2�tG��!wa�����5���y2D�s` M����(��E��r�p������5�"���
F���[�)}Ĉm�p.xp�8c�X�'�h#�/$�3����=��=P0u��w�M��s<���<BĦ��ͧj>'�&���.��vfY��ؚ�\�Ӗ�G`�(\��܇Z��,�A�&�!�T�G�&L��n���1��<��,c��ҮZ���pD�̲���a沾�jg��ͽ%;��r�%���'3�^|r����ַ���.���U�n)}��?l��J���ڲtY�t���7���J�������A��"$��D�|�)����p��vJ��?�����i��r�^5��a�=�V�_Q���츠R�V�톝����a ����Р�-�Â{8�K+V2�}��pPa�}����d�����T�<Ϻ���m�[����XdF�����S'�^���s�g^�k�^/�(�J��}JQ��du�];�as'g���� ������
)�<�#	I}'"S�x� G���%`HrS��5�(z?a���?��DP�J�?��gi�������C_��u<�r��~�3�O�?�;�h����Q�z�}�U����m��h4:�F�r�@�Aw��7��
�(F�p�M��6)�5%��A�~�d�r�+�uܟ�^(�#R/"�jWth9�L.��EQ}6�
����mM�1Bť ��ڴ�L��a�@�l��Y��y�#�A[�Ώ�a^���+T�1�BmF�n:΅+b�z�l�-�:&gp��y��w#{��A�Y,b��]��M9=����0�l���u���{�X��\��6-���"�`/����"����}̅]�]旰g����) �Jʻ���̌�։�S�H�rgO��=C��|�l�c6�/>'b{����jL�6���E(5��CH��(����5���h��yww��|��@a��î�D��|�+��� �EA���IBO�;�hzh�)J�?��D����Tac=
�1r�m�i�)	��:��!}^��}����q,�i,Jי�$nzI&���~貋�-�M�_'U�Zu���<��V˨����Aմ�ܳx�%�o$u�*;d�{�ށ.��l�Lh�$W?'{��}|İ����t�\պ�Zo�
�	�����S"df��/G=G8HV�L���%.�cTJB���7ja��{�D?yz�"����T+�L& �A���U/���؂�A�qU�'T���n��i����� 3}6��2�9��n��%���<�3tsL����/����ʫ�9�g�%j�G�:;�3 �������:��Bz.D��H]��qn}�8!ܝ ?O��yICߩ;�?�rѬ��^7P��H�������U�����oy���h����s��"]Mg�5?=)W�Z񟺣��_�x!��=4n~�����,�*Q�K����g%�"�u�ڔ���匝t�ߨ%Q杅7��@OzSg�~�#i+ʸd�8B�U&�X�H(����e����� ��ٚd�8�f�ҭ�pT��OX �4e����������U�0~"�'c��
@���	֙K&�')���*�Ԕ������_H@��Y[s�#�O�M���<�tw}�E�05��P�|���X��W��<�~��P�Ŷ��<���Hr��Q�Q��wM��״����o^��{]���B,�'Md�%h(e���Kh����]�̀�	��A,FolO-5r�-�?�&GF�'>��a���R)����Y�X3����x�$DO^.Z�2��9�VW�+Z��4O���m7����{����`��K�l/j��X�YGՠ� �p�N(�#��dl^���Y��~⹟6}��+P��%�0HG�}H4�R�@�R�P�ƺ2�|!�)J�uk~���p��}a$��f[M�*.8M?��rΫ��g�G_z��(jP��ʀ��#� �1�߰ld>��ۑ�a�|+>n�M����N�eI�n�9�=
�p�mv>�ec3�~.�PU��>d�B+��v ��?�e�u%��}3��ě�4 ��cFA����Zܠ7���J��H��gu�;?����h�� 髚z������A���oA����h,\=^�5�K���@	��X+�':�"s^b!d��?9*��Y�^�72�^��79�1<��3�G�'s"��"O���%I>c�7/�s��@g\ݬ��O���C%wU�~�m�Oקl�
���eI�bB�3�JȻ�&:~k&{Mr�R�F�B�Sg���"��l^o��&�'SgH�M�/�z��J����Y�,����px����=��WeP�D�i�+	�#&t=rn����}����.
b�v�,�h����m�;*$p�Nկ�5�@�`o��]���l�وխ�.U=���G7NУ����,�]�O��h����OK\�=}���ۣ�L�5т�����O��ɠ�[��cF�^9�Ǫ*?�Pz^�ne��su���O�n{���Ǘ��S9�啕��w��.�{d�Zc��f]F0+x���e���6����U��Ӗ5� �'��f%"蓂��ʿ�����������%,>kF�˽�̅9)w�:���fF�Me
$���8i�T���Ѐw�B�\��:��p>�-7-(+����}-���@��'5�������{d��a=��w�
�*�~s��Le�;��9Jg�d7��q`�@fr�4�¿�f���|��3�2�ˣ�)?>�Q�ic@����5u�({8v��,���UR�qt����(JjTع���ƗȎ	;k�p�v��*B<d�$I�S�^?ܰ̓N
�j���3j�L9�fx��YE�A$&��I>x���U��dNx�)�K.�� �����=�[m��>�q�O.����B�LOr��}^YB�:�{l�����#���*5n�g��H�rb��8;�N��^��(7��NEJ�ē�~�a��V��r��ȸ�T*�.��N���P���;��@*9��޻��נ����a���k^`�dG����C۵�l�Ŵ")���ܩ�����H]�P�����ah���@a-g.5��y.� ���qN<��xZ��O�k?���M!a-@�F�	V�����B�u�:vnA�m�ӢD^Ý�����o��&{4{��z$��_MX!D?��q@��Pz��Me*q"P�����<�m�j��Almm��0��P�T�	d��j�a�EXtH1F�|�z�zoʹa|A�C� H�V�؃)�_����S1�'��`�'�=���d�MI���*���t��09��-�
f�ptΕ�KJ?>�w遚�Z��.��G�vpv�h+����u�s
iT��txڋ�	�x���������,_J� Wġ�-�V9>���¬n	���8$f{�щی�H���#�@��:�����G�S��glD
�0�:�4y����I�,f�YE�wu�� ǖ�n�1�#��v�hq��b�%�%m��xg�$ENȦ ,�|�!���4a����S�U`�~so��/
]�H(!�wVh~qx��OU���\�?��:�N0�42�f/��¤�{FD�ǽ������{ц�5OXNBs�a>(� P^(��P ÜBQ�����ѝ���B���xJ���P�e�����7Q�NF�zěV�� ���!"~�n�A�2�^2�K���P-?.�	g�N��yس��,��v�p��e���N��=� l���gy)~vm&�_ʖi��D4��II�g�/6iG"�І��HЇ�c�� ��N���fh���T�`	l�xN�U�b"�O�9�v)�ʥ}��Qf)g<n�l⌠�S����N���DT�ǩ���m:�;��ݨ)�m��31a ����M��Q)	�����>{a�s�%Պ'��o M���+��׶q��(���\H�ahҔ7��)�n�>�ne����`�1z#pJ3��b�ǈG��?"�CZ��[q�"�*�,����O��;
��}�y^��K��//���T�gEֿ[�zP�O�c���̰��E��gf���d�(����˙_x��͙�=Y�9L�X���r��)�Ya�Hi��Ɂ+il���hڑNx|"|���H���B��Q�w���[��Հ]��cG�Z/$j��H�Wn�:�vf��/5�d��貞S��z{��q�kt����R \d���5#K�v>\�������룒?7<=��5o+VP�ڂ|���5�	�̕1�U/�N����J���V&��۹�`�夤L_��N'a��Z-�^�}>`��3�f����Cdsz��|�%��{�ސX��2�{Ǎ�;����"��xA�fXco��o�RAW��b�RY%�!�鷙0������-�Q��t�n����r���I &C�b�h������z �F7��C29��ʚ$�yI��5aҁ�Gok%��I;�):0:6��rf> �����+N|H����o���������MCr��kj�Yg�2�z����e͖�).�������f��K�L^ ����=�h}-���ذ����=��C�m��M%%�f(�ν����%
fa?�KE�`�)�bm�z��z�$��E��g����(5.�L5A&�*;�f�"�k�������:j��&�֞�:B�"1yˑ��XRWM���jkT��[t�ܸ�������i��@��EN��:Z���挶G�f)�N=�Y���ROC����9-4�l���-1\J�n�::�gE�����`��[�!3�I�c�5�Y#I�/��B��� ��e������A�&��j�����3LW6L#e�Ԩm\z+��y��z��k[;?�� �Iq���Y��?$8~�/�|1M�gԢ�<��gZ�Z�Qh;�j��X*R�T��� W�s���B�ބ��~t�\H�$��ęp�qi%��YT�Ɉ� �_�+ ��"9�N�{��[ �qsx�2��&�K(�i�]$���|G��Q���o�<G�w��)*�h�E����X�#��g��9�!,ί�S\�� �$��-b��ٳA�_�ʈ�S�Pe���MF ����^�|}R;n���ƅ/"�xx$P��Ň?Xf3/葬��Fo��+v�֨:�>
��V�6��&3$�����A�����cp�f a�f���hM�޴lYv.D['�n��\Y�2Ս9�0�#��6��	�L��8x��a�i��tJ��gq��r�Αh�nR�Å��	�;��-�t%a��U��G%�"��ް(`�;v�AO�X���3.�)��� ^�y]�I�ؙ�<���H"����}.kȪ�y;b"	����M�'�iL�sf՚Y���GB�h�p��L�P�|�xK���	��%��J
k_E� ��˂��
��}��5��]	��|wom��������7��IѾ���x�W���N������G(j�P��!�#�g�@M������lk�̇��
�K�O����ǣ��s�s�V�Ѿ[��dAJd&�!-��t.�&z�)SS���=t�׺}�U��D�/�t�E��R`��Q����9M>Dj� �gX?��7�����JE?��`&D)9�H��9U���Mq�9/�6�~�r��=`{l�p���CCc S�uqCX��1��m�c��v�A��W�\���d��&�n�j�D��˭��y�cM[��V�N�����(�(����+�$7�]����1��#<����c�;�:0�K㍬&�O@�2�l�&��X�&�ߎd'�e׈���Y�ڂbJں$�]�j��Y ��ǲ��|�Z�^���']�F4A�Eu�>��`l)��2������k)s��$s��U}�q�[�/���c�:Hb&D��ς�ZT�����ݺ �f*Os�WX�1�VΚ�?.�&#��So��,;5��ބק3eA3����0��o�]�k�rb�� C1$y@cĆ.>)	�M�V�Z�C����?Z�y"d �0C��la��������u'9�\�^z����
��9�M�D~j���hݯ�U���'�A�1�a�����k�������ɬ5F��
j�3n%�<�� j ���+�ԋ�E?O_	�T�8A۪]�� ��#�݂<� Q+�*�E[�40����!�E�	��@��^!��F<������<�]*�i��>����6-�*�=��$I֙�dvk�.���h��'�=�u��������^�\-_3���_] g�9��1)�h�cˏ-Q����wM�ӳ�փD�H��;$K"]�Jf>��V�#j��q����v�2Чa��7��;S%����1����	��s��%��tº[/껏��H�_������R�d�A[�՗��q�-�\̍���4���1