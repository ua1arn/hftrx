��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V���"WYj����i� �N�7A!�@<e�]ң�;��5DXL�%�����f�"|���\y�]d4�V���(h��_Ϣqn���RL�/� 8�OK���a�Z����IL܅T?5
�Nx0��Ϳ�7͋)]��2�� ���S-��<�&42OƱ�%�N�H�s��)}��Lo,����;��?��'[\�W_ ���������=��hm@W�)�c[~+�!?���Y�ƊJ�ΰy��Nh����ɘY�[�,�x8����Ί`Ա�W���=J��������%���/��>�Ť=5�+|���3zb�
�%,� ��)���o�ߧ�9H[55���	Z�^��u�_��Y�S�OJ��y;��18��"c�$���:#�E}�$�#oعV�Kl"�����������~ܝy��o���
z�o��[����Q�	,��<���"X�[80�X����*��@����N:atn<�1�@�A���#4:E�
�@��� �M��c����qs��>Y>>�_������
�|W-z]瓲I�W+E�N��H�=�w8���WF��Y�L�OH��͡ŷ�^���e��h�$Iv��Y#9 1A�Fl���_�}�#D%�����o~ۦ�(W�Ci����'�te\��0v,���EPT�qm(�n�^����?E����ɾ���wb����߬1�s>�:�E�d$(�� �%2��B<�-��n	2sSuHt������U�K�e�I#�C�i
WU*R6L:�z�<e��~�3�P�;�G������w�f��qAk�2PR@n	�Xടb9�g%��-���#��U,���7�����Ws��hd��i���;v��@��C
W�yi�Q���*��o/����*Q�}ry��V&3Z���a��O;uQ�@-�E�&��������}@�m�d����*�e�����ћ_����
����!�lI �&�*t�̅^aug�(�w�DAu�g�(섆I:Ũ�w���1�F����o9G�ٗ��ɔpy�ML�i����ǚ�ADV��J9��pl�<`�`�af�8�N���>�G�:�eG��N�^���2�"ל|�R�j��-8�E��n.(['g�7�<V<N�﯆��7M��f�c��?a���%D1��J�Q�^�)k|i
��r���q`�0�5Lz{���H_�T\�GB��Y�s���6�[��z	%h��
a�]�<�j�7�'���ݛ��>Υ�W�t�����S����|fZ��>H��V�
�L��|Zr����_�MTG�y���}�wr%o�$DF�p ������A�e+7����"ae`��1�;ӰT�6�G3��F���4�x�͵��j �u���^�'�<��z<�6�Q���o��`޳�a�ч	�A�2%]�o��c^}l��A�mH:�O���,�l�9��_��Qte:ϭ]r����4��)��ג��"�2"�����v�.r$�a�.����#����Ϩ����A�7�+Lf�me�5gm,S��c���ȉ00��LM������L��b�|��������*���_�~�ƙ�y��l���B��P?Zz&с����Sϣ\Xk��A�3���G  �Rw��K���N��+�$\w��c�l�5�"pp;Z��h�]>�;@��0�m3�`�T�����*u�(ih�p+ )>�.�0�}�����x�8~�gP�"/`$�Ϙ)����b��! ���T�"��W#N��	R�{��c��N���/��\N�Thy�0�	6��LWfߦ��S+#,�K3���8��_�`�@AS�K'���>�����^��W�|����)~`[�jGgA9Zm	�y��9�Y_\�,'*�P�!�5r�CB�@�ٔX��޿�[�����@{�:�4� iʎ܋��:<Ұb?'�{qb-vg*K>L܋S�jl�z�e ��!�y�A�~6��l�ͅ����4�@xG?E���b����[s�Q��v)��*�CV7�,HZ(�+`��q��|�<�*��0�	3���Mԣ}�	���l7�k�~Yɒ��@�q��'������� ��Ȕ�F�&���Q7�p��iWV�1ן�u[8Gh��G���a�;|b�����d�@w.֘�P��|Ѡ�7\�Muw4�\@�?�0դ+
D�\6mH�Cl�*;Ĝ�x�ʧ�4��t���C%K�{�ПR�R�ɨt9���ŋ�;;'��2|b�)���!�wK��v��P�Z���٢ŒM��G��U�Kꁧ�?��:�®brJF"K����f����sJ���4p0��Y��-W;o�b���eD��0�}(<��A�_ȇ�"+�m�y|���~�׬��@�T�"�D��Qq����Q�9Q���ĵT{�D���������]��O@�����Ff��� ��x(��8w�T�HS�,?T2/\L��ۄ��`��!π����n�;�-[��$�X�YG�eJx��+�]��Dk�ω:Ȗ؅#ƫ�N+���S���_"%{C�	����t��B�x�X5T"��~��Y�ڧ#�T�Z	��O��S����耑`ٺ�Rj�¢��d��,�F��`�{�9�|��v�O�F���Gp�����³f'�^8 ��a��	��܁A}��:�Rowƅ�d���&�g���*M�8��:���Y���'d&NO�D���K����ˢ��+(�`�>z�I=RL���f�������r3�]T�3����pk���uZ��Z��\P��*��v�������k톪�
���U*�7 �ە������1��Α�����6�z$*FTg~�S�w��%5��!�#^n���lM��'w��gs8-J*������fN9���5���s�ډ���ќ�+Ȑ��ɀ5d(�s�Y�~(�V[s�Y�l�~�ݦ;�v_��1넾V[�~��H�01��ē]�d!>0uEp]<���E�g��f�IX����T3��~�1�a��}���cq4�����6m2�Y/�l��~zFQT��A5'���j���4B�&�y�f���20��r�j�m�<΀y�&45C�в��r� �B�4�F��B\��SC�O
�Yƙ�>7`��WT?A��wZ`Q�l$�a
��[, =Ć��$�+�7��y}��n@�s��H�h��	 �K�y0]�ïȲ@����8�֘��j��8��W=�N!$wk4�V���Чr�\}	�F��4�c��v�{]B�9��d�k�Kp
@�S�{�t}���f����7��c��K�� ,]=��Z��$t��]�rk&��*g�X}p�$:5�9�U���ڻ�L����F�3C*�U��$�+>�/��l������\}~������_[�WK�-�%�=B�*y��;9����ԅ\���Z��K�-b��zyK��h�*����Ī�6�Ƃ±v`q%�f�|kg�Z��#
�1�2<���=j��ɡ�K�*R�\����$ccŐ���Y>���<!۱��?W����SXY�ޯ�6�oM�x�|�!�T/�S�5�3�j��2>����x�0/��W�Q!��x��_�k�|��������
^c�*�w���f8�&���%�m�;6�+�4x���ع�
At�K?~F#�L'���V:�`�L^%����Dd���p$n��%�;�W�S���@���	��WV<s)���S���,Q\4
E�R4	��ӌj5��\Zh��i*�q-�o��-8۠N���b������N�z�B�����K�`pÚ�d��;��b�"T/}0��a~m�<aB� FU�!s�#�hh%Egl�}^���U�qЇ�WP��Z���U��.�����)��xe�v��`�0Ǧ.�b���_<���>sN�QS�+�s`�ɩ���8.���6�ϙ'�\���E6LnK	�����M�~ᯈ�	"�u��x����z҆Äm-;��-�}(�����w��/�[�S�Q���ܼ�%F��L�.���̵7O~���(�O�8��2,r������H��6gd��/�i��]�r�����D�cit.�)x�(^j���ѱ~bed����)�KX�g!h��E����	k�L�����|��5�����WV�k���qG�F"�+-�<h���X>�oѹ�/��O�ܴ����S}6