��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^��M�ԇ���z��$��;U��ū���{���>zIQ�t�����P�ܹ��\�+�վ�<y���ݨ.B��Ϲ9e�%+��m�.���eտ[s�b�EL8g�˪��C����1n<�Т���j�k�U�|i��3��=%,�@����z��43ZӽIYW<�� 2c;.�RT!�*+�t=�Ϩ^�U][�"�#�$`g�Vg+�~�2���,��kti�Y�}�z���D���m�A�YTs6[S�T�k�!F�����U�'f�9 �/B�4�;�['R�Ź���yl�E� XO�1@~��/so�
y��F.���4�<��`N��K]�"�g=��&�������}v���	�#F���dP���
��k�/�����h��'�F��X"�Cd�x���~*��ЮNGϯ�#LX4=g�G0F;^Q �(o"���6]	w|*p�Z_*�,�wp��s��k�R4��xrǄ@��� f�Q9��5$M``�̯�s͂N�˕4���l�#���ժ���/C�ɡ�S
ѿO}���H�hP�w�e�9��V�-#�����4��a��Z���.�R����(�ywuD�U��7�V]�ml����|���מ�����v#�]D9��#h��PmL+�_����[;(u���}ւ�Ѐ��/xF�A��&=���(^p�I)f-�A�~�4������	��\V����/4*g�4ߠm��d��*8������}k]�dQ�߭���OmPvLr�ےQ(�0l�"XDx0n9���F�T�#������~�%]�Tz�����n���Y�fM6|���ܷ&Y���D�{6ԅ�&����<hE����D��2�����1`��Y��ΗB��-u_+��Hy`�����q�<�<z��oY�4~y�|.���`1r�tVK��V�2�1�L:��=�VWJ>&x�ʍ{#~�c&R�x�%���:�=�e�p�u�Z��~V*��L-�p�g�����  U+�W���M�[����_a� �z�#�j5az�쯡�N�*��#�r�D��r.�}�'��D+�YCx��5�|��i�����9�z�~�wз�xpr�'J$�~#��
t�X@�)��l �=P�^����ՕeEoꪨ�'��D� ��<�I� �&����n��������^����x@�i� /ƾ��Y�a��12sv���嚘�^H�x���ʵt;;��!p�� �k�,��bU���@�Q��J,� �<��r¼D��!��_�X�x��' �Z�4b]���==���u9��iK_XԴz�-�(�S���� ~݄�J��T���hA��//,0�W� _���"X
	,u�wƕ�UD+A��joL�Rw��ӥ}Ʌ�S��7 ֡s0�cWѰ�?���a'G�.vo����
n+��o�ה|i��e{2��P����QE�	e�(�@�i�������~a$�E h�-X�-��f��Ӷf<�V�4Z	���#��G�y�l�Hu��aup�o֯�*�lb�λ(#@M��$�	�����*�7�g� -pp�2��2�~�.�e�$$���$�:����dy�3zݴ8U���2K�OO��i��[ݣ�̦�7����c]eA˭d^����b�08U�p	�÷IdGxm��v�ה�fN%�Nk� l۵]u���EV���ƜYaF��ݸ<8k��z�&*�Zҿ���4Z� 3�jV�Zh��F�:��>����4L���z��Ғ\/֮�wV������q���޸ҟT��F����~���u�Ƣ��Ml�=E��_Y�K�ۻ��	E��r���E4C��-��I�(��,�bҦ�G� ��o%��t*_z����R����#�z�p(�Xlb�Ye��s�;�=jU�o��>�6�jgぉg��<��r�8�|��b.0UV��T��.�Rᨛ��=ȑ�s���= �{j��zUӓ��B��@����~�w.Ɵ���"���l*�4a[�ūa����>5$�>#�r�MZ������	��V��·��<���㟄��i5#Mcr|�{=�߾@���a��@ڼ�o�����5��^$��,��OS����X0���yln�b�\&�=!.���IX�7pF��p`2�a29E�h�K��d!��O��7�o%ă���#�W�Áh��-Oh��T7��<?��-��Hs�*}+��wy��HʀAFl��i�"��tI��� �0#w�D���~�ޱ/��O��>Fm� tT�0����R�YR�B����3�����g�Y6�(�I�?o��.��r���H�ʐd�"�Ʊ�P��K�V��	��JOY}0yP��wi�>���Oz	MFǋл�P��卩�C:	��5z� �q�����ǁ��mA��� If�)�^����Ai�9��%6O!lN.Y�.ȗ2�fxwL��1�n'�����T�@r>:Y[·%�LA謈�Z!���t�������ʊ#�c�Cje����>�:�����{u���/V��}��P���|��P)~�6&�����}w/��oY�)a��lM����>�ڀ�z��O
2.$9��ߟ�L4;�V�H����r�ɬ�B����<��l\�O�lW̵�E{0�w����ڧ'��Bht X��͐ˇ�"6x�����[	�B��~_�	����dO(��ch��Ơ2���\�Ry�d;%��dM�^�u�A��M5
������2J�tI�Ջ�{E���়�L	P,�8�x��G����?`h_έ���,�a����f��&v�U�1�n]п2�/��=%�n�_/K�Q_�tHb��1�m-A	>+�l�a���O�')��h�d#��$6B�^�N�~�6Y�X�k�G!5&���l9���N�a�/���RB�!M �"7
��1���l�����"�w����P��*5�2����g��pP��7���G�8�1o����/�lNXQ)��f�&:k$��*����_X�6%U4�TK��?*�}����x<��:�"�Ҁ:3���b�dI2�GqQ,g�*ԗ�!]3U��HB�j��>Xk!���g���	����}��m���C���I̤�l�%��l����� ���,�1���m�5���|s��2�qa{ߴR7��FI)e�_�g!�e@&`�D���8���[����Y�P�&bF	ag
�u�l48�cX�h����0�D��	>q)C�R��!�ү\�p�a��g��۫�|�#R��-BV /���g�=�k��}�� Lom���ӫCR�9l%B��t،M�s��d��``U�6z)C�_!��� �d&�Y"����|m+k]��~l8�e.X2�V�.%0��<��$�L��=�X����Vp��!Z�QGm;�t�Ud3�s}�%�ଅb��03Ka�Տ����<LZ�aͣ�������`�ZGXjz]�y�)>gn~/C�v�/������ -5���� �L��� YU�i��X�RX���$Y��I@��q�8Y���}@Mr�L�8��mp$��VB0�P�H�PW5ґr��A캮n-��A7G�TQ� T\e|Dy�q�2��7~����*`j�q{���Kha�F�DF`��=h�	qC4�͛�@���aph*�������Ns��Zi1E��>�V'�w�:V�/Tƅ��E�[k����.|��#I~�IQ���ˀ8��3����5�x��,��b�F�!b�k{6����t��:lw���s�4�	�2[2F�/�fE�' �
٨�F�z��e��ږsF�0�������%�Ax#��W��eE��߱��&������]���Y�F�`0��v���H���*�kp��ߵ�!�#�`U6�H?��k����+c�-�t��V�֪�;��r=�U�<��6A��,�_�zc|Wq�����_֗v��,nT&ViaC˰�΋���a�g��H��j�3��$yŚT'ld`�K}7ޙ����	���.�?�7�HCt�'�6�8G�����T�ێKݔ�,JU�_��K�;���k'j>+�@\���o�Q�c��������qUz$�R�j{�͆"g"���P8�^�?a��ɛF-eNG�ħ��U�js>�2��u��~�*sQE-����zK�,,��7�2��9$�ؽ��;�3]o�D�rsA��o�X7]p|,�����AfJ��h
�҉��&��ᜒ�6��6���3�/	֗�S!����18�Bq��Β�е (vM�p%�5����5�0h!�8���|�Q�������[�]�J����	�N\�Z���8�-�P���.�xl��H��P��T�0�ځd��w�O���E�c~�+yFwV���o�ΐ��.��:�l��^OuE,������m���M�o�<az+l&�����@7ē�o�Q	�N�p�ݩ�#�I���7���O���5�є�6qX�� 6��F;���Hj�U���c�/ه��`-�h�]8�+��d&��ݺG'��bg��4]*1���_ʼ~r�3!Gql�~���z�ӟ=�Ww۬�W�'��/�U��tD����I�xP]nl�<;+�d���#��׫�8�{��ϕ�&��ׁ���:&on��4^'/[�s�+b;t.�5���*���;1<�
W0P�>��WH�*P�_��[�5�!$�Ƃ��[�Ȱ*��93bę�Yxc;.2���i3��dݩ3yJ�n��؇I�JE}ٛ��\ԥF _U�1/�f?�
�A����w�5�W�$�E�#�s�\���M�r�g�	�ФT�&V�n�n|��'���������n����^��z[]���t��%Xt���-�J_%ÓsyYU�(8�JV@�����k�ir���xB�p=fT,����Nx�����̖��7��E�����S�K^(�OL5��g9a�-�p�d�	K�)G�xy�]r�pG�����PbQgw�d���9�L�2���#Mb�X��l��>�ߑ�z�\��5ܗo�ifS7:�Q{��y�mP�	��Rz��}�"���t�i=���υO��ggC�2���ek��Kމ�ns�t���A��2NG]����؜�d��*�x:�<�\Y@p��8MU8Vo�м���U֊?m�k=w�p�+q2��\�p���Tǆ?%?[К3����FM0� 0�X^H��LO�4D&9t����Ӎa�h@���u�� EZ�0�Z5q@�9׬��m��e2/�MK��S��FE|��9���A�N ���h�鼂N����k��9�qF��8��Z���qj,G��Dnp�p�Z�࠺�9��Mh�R�j�H�����T�q��V��E����Z:���3I�A�	�/�<}2}�K�g�4�����*C�c퍄P���p��1(Hpqd����~�'҉|g�t4O'K|'B~�cGu��) � G;މ@ra~:�ib`��G#8q񫚸8Yڻ��ʐV���)�U�tg���,�K'}�@�BX$+β��cH~��~��^bBgTH,`S��$��яL�tZo����BV�?��5�ѿ���%�5�CN�T�^�R�,l�Ԙ�����H`�S����r
���t1E�U"
rxT �RfxdDK�3Pa����m��9m��n�p���g�`S����n,v��;<�S,ϠgQ�h�D���#i0$5t���!_�G��-�Qo����;�Ƕvk>`���Y}��V/�N?���
�L��'��lx�,�迭�h8���]���	膃e���1
^鲰5�rxU��] �űU3悩n��6"�xr�
�����3�<۟�;�-�E_���,M��������V�L��@�PMF�̓g�+,>?�(B�(���d����>H�_u��@�|�qUi�+\�d����Х���SK��q��?'��p&Tdu�Ժ��#�@�	�e�zԔ��5��_�)m&E�2�ƛ�㤚F�9XKd��Fm�#�޾�z�.q]��ڲ��a���T��=M�is�x{���eM�&���~��Ϟ���կQ�G�����7n��ʱ�d;�ڇs5�w�����:7����Wz��t[��H�������W�����))��C	�C���ԭ}0�Hۚ��BmK�Y�K�c����=��c��=XH�9�������ku�����Ό0N?��0�`�m�� M#n�mg3�oE����i�����3���}[Hs���K5���P�j4���k�9'>��(�)m��kg5�ȁ���=�fK�K�%%�((�P<j�I���Q��2�:ε�G� g$�A�Z�J(67:3-W�~���R	�i\4L�$�)��_S�>f�z�� ��;z*F�E������hJF�[� <�A�g��m0�4���~M�T�s�� d���>5�S)fB�hz�WǏx]����j���3�O^�����K@��C��si�������Ɏ���lY�BÕ���5�J�L1��Q
*�0�Rt����<a�Op��Ca`h�����o���-е�!˵�6�;uͲ��)�i˶:j��e�J�!`���]U��kr�6��b��a9`��bab��{�����(�8Xɗz?,U�$�Y^������z�/�h�G�����4��O��zw�ݝ9����u9���E��BshSI���F9��IfX�f�����_��\�ɸ���a@	o\�r�[�L6Ÿ{� z���H���֨�9���X�;7(=ĸ��b�m���a����PCַ�&�,�٭k��y�X8"�k��Zhl���8��Ё2{G�u�{}�����)������;�V��D0��A#iE�md!�Q��
��)������1ߋw}�ܿ�;���L�S}���]	�+4���)��5Ώ�r�Q��b���i?��V�&�7����h����#R��X�ve�� %���Q4u�ή� ��ҡ.���k���[�Ho�D����^2e����y�v��f�G�@�سN�0�Ι&��P	U_�t{A I�iu�����j73yB�FqU��&�����eo�9�����B�U58D�Y\K9MO"�L��W�2�So��S�E)B�ryk&8�Տ���xT�m�60a�q��F8�XA�D���[��;ɺ����R��<Ht0z-0쟨��]���E���y��Aas|����^4��~��eL�aןi\�6�RT%?-t8��݉9��U8}d�k�e���_�	�Ȇ�
��r�����:�k��6���$��Pd�}��G�J��y�mS�~�Q��g�㐜P@N���V��|���?Z���¶���#�(D��#W[#�X5�þb�F-��3/���3?�Z+�(a?�rP�p(�_!���~���X�d#�\�@�7�f��J�osL�I�s𮖜V6��y�ʴ:	|6 (�o\,N��=3��(�Ӹr��R6���G�8x B{��q�<W�p���<�L�B��=�I���3�>��z��t�2#��H~��i`F�w��̵	�l�A�+����;�Ղ�r�*a�zǯ]�fZph��q��2`/k�C���Q;Vg�{�Y?(�a��G�`�N���&Cs6.o�{@� �:)��ww	iի��J?;�g~>G��=Y/X��J����x�FHN*�K6ի%Z+^"�bC�SG��nx���6/��ז�
����&
�x5�|ο^=8`�����y^2f���Ba�N��ErQW?�56�9b�T||g������*��:}ђy���a��
*ñkke�ߖ��*QM��W�\5dO���D�72e�]@���@Ԝ���d�A�'��M@p�
;r���;�Y�j�[`aEO��ǒ�Q:��*u�񥍃/�jl�����2� ����W��H��4!͟�T�K��d�X�Oһ�Z��{�7��6���=A��<�<�CÅ^��\���� ���<�O:�
����p���?X����5NH�;*d�"c���R���,�)~ְH��T��6�,]Z�Ɓ�F��ڨ�N�������[-͟*���E�[T�}����v��h�+�� ��P���='KQ�H9�郘��#�|��P<��zX�k��	Y�}Ox��Ө�>��J�'�|�.Jy��Dg��A�Y���=t��뀷f��Y� ����=m��ܦg���J	�ڻ>۴����g�ߺ+ȏ^'�s'5�!k�8ٮ���|:*uT)zMfb_�q�Ђ��8P�)��4�z]�@x��B�@�^^SY[mkfF��b�n��c���Ӿ�z����"����IZ��N�L�L+���4r��Yp߫��F�v�(��Ӥ��3�B��{ⳈD�����Yp�j2�{՜k��}F�~$eԜgA���.W�
Y��5��c��	E�/U����`��
W�0�Hl���{�`qY�vd߀+�f�ʎO�（�	:�ȩbEh�]c�e�7.���[�]�4Z�A ���e5e~3>���l�`��;	��}T�ҁ�n��1%�pX;�,���X���+��l��'4}{�����Q�$j���쀇���cr�r(���W�W
鳨@>!�?	��H����>	�s�d��ER3�F`�#�|O��g;g�o�M�u`��پ=�r�x����6v�$��=y�+���$<�=��6Do���\�����~�.yy��e��W�]1�;!V�\���,>���.���@`��YM/�i�)�@}E^�-�`�ܺuo�v���s�@i�{p���B H�2R��d�>-����YN�y�8�h�V�~���[��6n'ǫ�$�CK,�qr����K��͑��ūWd��+��|o����o�u��LK힭�n�^��F�ջ|�A=)��1�JW�gyn�]���1�V�$a�q%¹C�q���I ��B����� ��M��a�����$�����>B?)�N��E,$���d��@�������T�B�RP�� \v�i_�/��!fBU"cC[9' ]��$�ቋ=AW[4�G���GC6���䜽�wG��U��\*x=�)���T�a*&��`�|K*�y}%w'�u%��}k�.� 7_>�|"��1���c} �H��L�rY��U�<Yjy����;���א@���F��lOE$��q��G���kHU��r��%�f�4:�P�Wq����M�s[<>!�ґf��B��&��i0U�:�^�)k�l��_'��4����p�Y�c�����l�ċg���jz�.�+U���q���T���5맮0�{GȻ�P[Ό넥h7���Z.�~��F�B��^���� �v}���_*�Ʉx��0O�v��ycf����2��E��R�[F��구���"�r�>�=Lr;�/�r&�/g��3u�Yn&i�a�ﷺ$�)��k���x�A��Es_-
Z�8�E�.3���E{m"�y:Ts/�h-4V'������~�lR�
%�ғ+�`v�r���� d_����k����`�9~���}���$t�������`�E���#:�!/T�x�(ϒ�,K�F��7<Z�LZYy���6Dd����W+�6�X�	xAq� �g��e�P$]�0�֢���u+�j#F���i?zW��_L^��u}�q"H��������$�q���"���#�#�?
��7p�۠�����[[%���q�@'-L�uu+���n�>+��@*1�@^-&^�
ɐ���bn8j� "W�7��Z���J��F��.+��g��9;�V�]jd� K�n9�����x�%�_�!K�\���n��T��
�V�š�{7av�!2~���R4� ��ե��U�P����Hә*�zӆkA�p�z%�"J��7�T	.�ZdژW��ݙ�qr�d��}d|��̞�d��z�� ��u��?�wXX���wR�A����(N�k�E��W�1���n����z�� �m�b.�!.&�]_�l�p���d^�����|���ZW�_��M>��7�%��7ZWw)���Y����Gv;]G���o��Y#�`�_�:鷉����޶�<<���~W3u��V�%M��A˩�}��C�!�mY���@N\ T�D�`X�Irj7�*V�N�_��^+NBu�A-GO����ہ��x��0]�r��p7�Ⱥ}⢁��+rO𐫛�k���h߁�5}����8,tFF�f����'[��hdLAp��k�} (��l}��K+�iȎ<l�W���5T������|{��Tp�0���@*k��"tg�#e8!|�n�DK��=;��jہ�p( yoՓ�.�v%RD1�q�	�`U�����X�p"s�j�J�>;�<�Ģp�u�Q�!=��1T;9l�\Z�g.)��(2�yJ�lhG������={$����Y��o������p��݈�ޒf0Z��w:u��\���q�A-�v)�(է�.To����f��� ��
�_,��h�k,� �}�}g������Dp�z�n�<Z\��1����0.pJ� n�Y�2'R��.��?���̂���G����BС��^ې�1�4��'��[I�ݯbM�7�QHV����=���bM �I��/�� ����E[��&6J�S��o�'W9�K��vCs7@�4S��3�p5��WLu��b�j�ɂ�V�0[Ф���+�� �V7��4T9ul��<[||v��l���-�ͽZ���2/+"+,Gf�*�)�Y6��X�R �^�~,ϾuG3sc����$�ެ}2dB^	��хh^�/5�"[mB��C+�$�)�����J0)��|��1M���h&��S$�IHE�r2k�L��I�/aS��	,���jnp $d7*n��J��E��V�f+�W�QG��7g,
�a���RS[�>}��~�0Ps���op)�$K�q[zz$3�4��#1�����ο�!��9-�r����V���I m1x�{��c�x�r��R�;�a��3V� �\����� �[�r�"�����	|�^���Ǫυ-c�G��Y��K��t�{�ěh�w�F�bV;�Y}h��L\_���q���8kF$��\���#�D�V�*�:��b�rf@�0����=�;��̞�;��!��0�gr���!5٢���!d����;8}����Of���F>yw�%��\������֏��FdU&�Ω�G;��� ��U���1_0x�6C١�ş�G�������>b�=�}���󭥘u�l�h&;�,[���,��S�u���;̭���2
���[r���:W��3	F�D9����=���[�����;$&����Nd�a����N�0�毐���>������G {�$�	�ܥ�#�LT_uF�z�#���~em�\Ub-�}���W[�j�V{��<�:�T}ȹ��7Y��u8�R��7%�p5�(�nzt�~�R)N�}��.�>�J{�x@^�_��^�ˠ�D)��Ja�i�Z�^�i������`5�Vvy�G��E��yݰ7�F*-��٩Ӟ�ۑbI��k�8V? L
l�1q
L)�cK���o��LxB��
s�x[�DZ����{���W���ӻ���AA��5T[��q<�Ug_l�9�HS������|����?D���jj���ȜjW�
�~�L�rS��3�F�_���ٿl\�ofB��(��Pa���G�|��؁'}��G��u�����bS'
���,�M
��L]W`f�������d�°+�^7�v���-�� ��OQ,�;��kI��9}�M�k�Μ�9����%*4磇H
,G�{�IE��&�c'��N�inu?��:6�]G^s�X�[�ڸTR_�����!��s�LU��1��4|��`�3�{�	����W���^�	��{��� �FD�_\4���3+�M��)W�(9���w=����Bq��y҃��6(�3�׫|%/�$�!���'j~[��Q��>�k<�
��{4�6EqY��[���m(��|��Ć����>�p&���E�����ο�ڒ�iwT
�?q�~�̝����!���&������q��4e�-�tŌ@@Oy�V�@����x���U�o��KO��tV��A:"KƔT������$��X�#�����k9}i�W�y�Y!t��|?�}D���g'��n��zӧ���E�nb^��N��-�J��v�ajX�ۤ2c��:M���4��}�W|Q��4;x���Ţh��u�<��H�6�_�(��ߑ]
�X���ډ������[�����D�ͣ�ދ4e�NR�$���RC�1��v���kP���H�o��;s��k����)�>&|�EQ��������������N�2�t8![Y$��tL6#�|�N�q���UHA���X�I�����7-�ա�T{ļŻ�7`�ԅ�����B�i(�o2[��DV�p�r\&}6���K�(Y�g&�@���R��r���O	�D_�-���<5[��L�39�%h�+��	��Dk�΋��y��)�PHV �wǏ�)��2}�N��oT�Ɲ�}�([N�F�盝�W�d��L�����稥`ۘ��Zm]Am�z����c�	)iTĉ�4	�v�\�F�JDD������v���<��j9�v�M(��O��t��[~��lv���_u$���	�����t6%�A��Q�J'jLn��S�0.3�2O��^1k9�j�VK|N�,����m���j�D%Y�sW���h���/ڰ4�^e1���@��?���� ���aA(�>��u#y�6�}l���b$�(�1��m��+�N�����G����V&[�@:�g������F=��$��������#x�����d�ǚ����F:Ӭ7�P6��{e�l���1X������ɚ�d��5w	0H�#*o2�-�9��0��ˎ�C����i��A����R_����/W��ROb��*����o�L<�wk�������]-�}�]�۞��ƅ��z�E�rˏ��$O'�*daOv�|c���f=$�{r���K�K��������w����M(�b�J�x�G��h��Lh�!Z:<��A1�W@��((�7q�q�T��:���� ճޯJ�]X�C�r����Ng��
f����˒ G�<?�1�p���f��(�Di'���@b�ʏm_߀���&=�}���^�InϚ�!ߺ�|Ѭ��A�0z��:�A�9<a��l�c��Ѹ���ihG��C	r�|8�}{#�+oq�a���h���{�PqI2]s�j�?�'����EM�{��F��X�6PJ���~��{��s��&|/�S��V��&�zR T0i��j�,<�qJ:q]>r��Ku�Wf��3l�?f�� �Pk�'��N=��}�LR۟�z7���sL"���V���t��4�i�:E�c,�����g�̊�����:
mF��>��>r'�blS�� ]h�c�:�k$&��}�S���pyQ�\H�T������{�)���rO��.0x)˞�MH�L12�a�
0�N7	��9c�U0�?����l��<��Ue����v��8eH�m�̓���.-
��0�>��&�`�#�v}�����l�V�pw�ޢ#���o�;�	n�Mr4�~�{��f7�_����;&���e)��W��_f.wQT,�h���Ȝ`	�gm�X�!�~L�P�f��C9h�	˔�uD"��K6ˋ�-z����;�ۡMm�+���
&��-�P}�o]��"r���Md�D�hf�������B�	"^i?a*��J��3�hq5���*g��_�6�(Z�0�f��o�#�k�Ck�������<(4��-�`�·�����x@�fCb�}P��6&�UTI��D����	H�$���-w���.KY�b�T�Eŧ���P���è`�U�k��ꇀ� ��c����ĽG��%��۸�{����b�D����_����o�+����jC=<�)�y:P"<��ƣpG��Ih�����
SB�ؙ%�fڎs|.&�B�����7��pW��*�#EĽ����{8a6wp=�}�OT��4���9sɥ�"#�٢�P��y)�'6����Ha��j\�)���DT	�~�B�>�,��t�e��̌0�BEk<mv��>�瓩�{�%�-�;,�jd�K��*��m�`9��4v�|U���e{.�d�����bG*R���)A��z[ŮG�\n��B���$)D�1���hɒ<���N����˯n/��h�� �y��D�=��5-��~E���N.����o6,���������&���)�Y�w�x�j4�{C:�?�ͭ��W�v�>�p 9۟����$L��ʶJ�O��MB�oUϖ�0l`GƂ�w
bGƞ�8�"���Ehz�Yۜy`�8�5�nj������ub�\z��񼣳[�b���;%J���{�瀑�� e$5��fL� �1$*��o uBh���jC���l�xO��8ζ�w{/,�0��rP�@�Q�&�k4;4�^�1P�:���̵�xc:�|�FW�6��!oU)j>�s��~aPR��.��M�:=Cnn��z8������ΰ�����(Sh��0�z]�t&|�c$Ҵq�%O�-�&&�RJ�P>Gy,~yʫw)���L��>�>P��q�2���+a�>��<"� ���������6WbVv���D�˘��R�yG�W���=�K��6o�?=�w?���ݽ����*Lh��k�&'���� �?���D�r����O�����:�ڰ��y�$9V@�Է����Ԉ�(����归��k��)Yֶ;�/<e'°�C�ΜA��(UOL���bψ(�#&8$�wp��V�{�>E�&g��;��6Կ�,�L��Y)�k5��6�2b��.4���ʒ�(F�r徨���*��uY��G���pN1�t�"�]1m�'(b��d��.�j������!�(ѥ��a$oR��#cU�����\������e���]��<+�Ce�A>�G�ٗc�J�4�TUe/�7�G�Q�͈�Nz��S�������c���;��Yf?w���ф����˕�/mxy΄%�X��"p��ʘx���$��a!>Bb�w���~�"Pb����ɏ ��s����\ܹ���o�NҺ��=�г��%S����� G�_��YX�f���h C�=h�jYʊ�+NL�_Z��0�FVU���r�R��86?|*��U�W{�r���ఈ٦��;��B�IRڏ�$ŎGç�p�Ն�:.��2��~��c�F����ڝ���s���_�q�A�����YK�+O�a��!��LI�:U���;�߾�d&�O����0�����8H�	~yoW)1�/��TJX:��n�yX�5��IoN&}������N�Q�9K}!�0��e�l���Q��8S���W�	�
����{�%�N+�"�N��J��L�eB��3p��� `�(���?9��-��L~h����rk̟���'1r�Tf�n�Ә���a?a!"Գw��+h�����	4m��a�>#fZ���j�:^�Pc��y.�����/נo�ƫZC6��^߇�����
Y� ���H
��~��%U4�E�(�Pr��CV�[�BO��u�<�����c��?8@����4�#��J&��[��8uY�1K������ %���#JD|��͓#�+bwI�)B4D��r���t�a��y.C:�����ݡcgq�^M8 &T/�א��C��E����S>��Y�%Bؠ��㲛���o�����K
P1��Y�'=�Z�� 1�4�!�VN!�Zb��'��="��:̘
�V����)+��]�C�t��<��s�A�f���=���#�R@��J���4cc�	���)M|�w�=-N��J��Z��E����k~|���U�b�`M�����`r��ʖD�s9{���u��_!�Io.1�:)o���f�R�:4\��>c�Wr�~�5T���Ra��b���C�A���ʍz����,���6�t:�/܎/��F�{�딘C�
����kЀn갣盩�����ע,�����k�_����;���x��6(`a���q��&�@�:=6��I�cm���K�KSe�H�T��[�&eb�螫I 11�;�r�T:<z6?�*Qo؜2�\%�k��E5Rv��G�����B%{��W��~N��ń{��Ԩ�M�nq��7��DO�w����:݌��Ӳ�l��e�n�E��㯵���snh�C
�'�r5�ڛo�b;J�qއhm? �P�nR�����͡��
�y=е\�K��e��,�JC��<F��W�$���`p(;j�v=�߉��lvq��Bw�}m�{Q��C��?�ckS��x��g���h�z������^6-�sTαn_�}�x�wQ����%��� ��+�:!�+Bc͇M�wB���ü�*V�Lu
�����#��lx�	�:��ݪ�\;ʠM�1�VX��&������!��b�3�#�y��,��T��;�^���M�j_c�i2�06�:�Ak���ԣݮ��	S|<���C#���v�,��m��W�'�዆�t3<Ne��B��%�I�)jv�=t�@�(�II�4�e��*z���xn�s���w���8dOmr����4�{>���&��]�bln�bP�X}؄SN�)�ܓ�ˠ&�U,�K��8Y��9F{����_k͵(a�i�V��Ŷ�ܖj�;N�q[Wd"��3��T���f��ۤ�KdvQ�c�@� ��Y��w�7xLq�5�� =\�0��Iڿ.��d���C@l��~�&ia���3#ڪ��Q \����m�u�@;�Hi�@ބ�M��]��$�Fݼ�j�ƤR��fЩ�t!c��s���v%Cu���.)f�|�,#]xb]���t�Y>@�H���iS��bQ��],(���h=9Qs�F�ը���^<���(N%US �"��G��T�l�B#�i�6c�}��㋒;�<�cyQ3�*}�xk���|�9?M�UH��b���V�T����H�7���X���n��sT��sBK)M�3Ak%Db�Ĕ��`k�5��|!�ܮ��oj��z8�����)��,|-��G��s��#�<�VzxŌT�V�?Y��mY^�M�ˏҶ)��,���о�VE �K �Xޖ�ԽO���p�nv�x����d�Fd]�S��'��}���.��[ _c��f�0��u<9%��Z�f��iKG����&>C�֢e[1c�t��p�<>9�k��5���P��\���
�me�iH��i)n'6��&�z�Ft|O-^CgW����Nv+�P^O���9<M�.�3u���@���u<&a"������P�B�'�����qE�9S;�ReX�[j�/�j&W���cSB���bԺi;5��[�Ӫ�8�|�
���ȉ,��R'6��l�9e�~�&δ��Cl�n��0������/�f��Na�+�2�q�Ӽ�T�j��ϊ�<@$F�,>�_D$y�GY��aY�@���ۯ�>����1C�s;ۆ�F2dq�T�h�5�3�ad�dĨ*G��B#@A��z'��~���B8IR�mE̵������,|`�%̞kz�pL����׌�$TbH�e�A�"x���F��-Њ�l�x�R���1�`�&x�ٓ6��w�XW�NI{�����0�=���8�a����I\�a�b�(�_��A�	�>���~��ֈ����BWβ��l���(�5:�9U-�;E�D�F{�g����'���ܞ�c��E�w�PN`����*.��t�ܴ(��?7����\)�<	T�_
�z`A�Z|���T4s nR'����iK �?�����gv��KR<i���� P�`7l�J�e��z�w��?�И�jXw�I�O�h��8���3��< 4r�H񼢗	-��:�%�[$~ g�+:���q�smnDt����q�8 �=?k�� ��sv���F��-�P��v�d/�bE(wכnW�E}�Z)TgdBg�]�l��S��]�Ќ�?��\��f�^x���el�6܍�y@����p�
)� �����xO��Iϱ��ӥ]i��H�٭uujLc�N�)��Xk-�ꗪ�!F���)��uث�i6�3�Z�9,�5Mא䒅F(αY��#��9��=!\�a�?��9���4�}B� 3O������NTվ��|5�ϳ������M�I[�Zΰ��bO^ч��}�&Q���z�V�궺Q��\o��M�N��x���}9�dh��Z9߲M��r:��(Ŕ����B��s��QQ���Q���}ϴ�U�<` �j�9�]Y�e�!�u��Rg�˒W���r�
4/S~�v��੣���4aJ]z�K���.��A�ǜ��w��<�V�7���Ŝ|l�`�W��%��Y���G1e��$C������	s^c ��Q�L���������Ƙj?#M-�?�,��D�v��u���fQ��Ǟ2���+�!�N�ѭ:?킁��ҝ>K�Nu�SRD�(Љ�~[�X�:K����?��	���B�l��pII�Au���v����؆5	��{����i�,5�,��'5�Zas7�ȕ�i�[F�4%Z�Y �Ip���6~��%P�c �-AjȪ�n���� ��L}?�;�q��Vb�<z���l���X�H_�V��Ց$�Nt`�;�k��C�z�7�4�D��.��0*MSgr��+���x��o��Y��_\�8p��J'M��H�� Ue[K�(/��Nn���;˦�z�wp�3u�Xp(Y�Lc<�A̘��x��h�HNOj �����=堟����.�|?P5�gp�B�R�`�D~��7������ɒ�d�x�E����s}bl���Fnғ���w{�v��	�uz�6�bQ��$�+(d^�gX4ȅ�	?�.��V�n�l�@�$����{.����<���4ۓP�o�e߮
��0i�p��w�te.�����x6Ot*��8��d�lҘ��>�Nz��ߑ�±PA��B%bmۭ���q�ӝ�J�:��8{��tHl֡��j�̭S��E��O|4��˴����c:V,��8C���� k�Ut`�v�GXcX���}�n��=r���y���M$�����Pef��"g59r���H�3_Q�٨b��z^g&9�C��޺�k꫰-��aK�G����'̢B����Ԫ�`R�ۗ��>�1Z~5&��Jv���a��9kA ϯiJߧl ��7��4�W/ڙْt]&|[v� �@Cn�T��	c�d#���-B��5h�}�%l�(���Z2|tb��eTE!�z�د��k6���\��b��C�3]��w�}򨴪<=�� �z���E��r��(���L&��[��٣$�]`ӷ%R�k؝�~^+'Y=�^	k���t�A���_���Â$!nT�B��ceє�F@����X�sO߱�U�{)wB�p�ތ��:���y��NT*5�䝥����~o�9�kD�Z�x����N�뎶�C��v9Qg��S��i�|��ߜ�)#�R�s
BFh�[�S�����ӻ�L2��>jΒX�l�9cf����8���8�܏�2���F��G��� I�*�7ݙ�B=����sC�qٵe�ֿ #6���؛+�X^ٕ��-̿�)����\A�֬�s�&����]��1q��,�sPg�Y�v�I"�B�&�:����_�vx�O3�1e5)G��nc�Ⱥ.A��>>j3��#L	���;n��7h's��Bҟ��ŝ���׋��п���W��5K?md�a�V�Z��ǟdr06]JY�;�D,��:_i�E0s��!�����,oL"��ӱe�:j�۽y�7�~��\t�61`XTh]�+{F�
<�I4H�u��H��B�8�i&o��[.�Q*���h��ţ0��ϾU�h�-#\@�T=�*���+喸��	e��c����0�U�A�(E���$
V��O���R��/���2�^`<����g�w���Ǚ��y2k���auͧ慯>^��?���?�ú����݂�
�D��U[[Lk7(kw~ �K	Ș���<6���Ll˸��� �ku4����_�l�c5�>|�g��Ս�g����B�U�t���F�O�I�1��h3N�I��7|,	�k�xi�@%O�S�<9?�Qв�`�����T�~�g�����?Q��F�S���z�d���!SޗF���抻I��Yc�Vn!��m�/�xt�"0�:�G%�����è���e.��=-�r<� w*!wl-e��\�\���h��8<�n���Kcޕ�C5��e�b��%�������5�Q?ҨWw��L�Him�^H��$�}�2�Se\,@��
v͂�Q�D<
�!~��}�:��dO�[(.&�@S渐$��΀�iu���s��*��0G��@�������M0��a�0&or+��%����e���w�	���Jӽf*P^��`��~tMl�r���xL7��xuz�Ɍv����S�G8j����E<�g��^f z23�JZ�!U����8mYЭ�J�z�b}�����3Q/�bI����	����2��AMA@����U{�`ȴ���q"�����Bk
�1�� &��R��͸dY�Ȕ�n4�,y�#2~(b�R �_�Q,s~!�=�"��觛u��<�^,0�x���43e�Lei="���{��3�H�]�ն9�=�d"%�J.�=�C�BLoJ ]]�Mc���]0��#�6�[�����6eSwK�:�(7O�]i2C��ʺVْX�����P����R`�͘5��롓�:(?t�	-��skD�1��s��rt�u^�	C'4���������_t$�H�_]P�*�e��C��:y���"N���^�Bvz!��I���ZxH��?/��jհ�7�&�1���w��P�(���VP�c���`�7W	?ҡ��Z��{��s��>���D��B���J�b3Q�0����wE3�C�S����z��E*�Qk�9�@�\��~��ʇv�@�jB����i���;L^�v���y��H-�֎����$��K܉rr�fÅ��<��3�lh-�$�����u	�2¢��T��:�����5��6��C����%���6:�v:���]�Xu���}{@���}<Z���d���j͊L+��DA�*��V 4%?�����P�@ن{bчu�+� >��<�a!��:�[te&��ϥ[�j���u�<=G��>���9#i�+gȈ��5��.C_ګQ���m�^-�s]��������@�����>`�=}qe��6vܞ��� UPe��,�s}fږ)(%CP���=-"}J��������&Pp�;�G�&?����n�$c����uC\�yz����]si��tJ���9�"I;���*,'���n�H�U�-7��xqJ�Ǎ{;�����3�/:�J�ѭ�r�Cm:�����*u�q��n��%�/��B����������TK�~V�=u�yTiN�6GH�_I:�j��n�	�����zF�+�'�3朷��2R�[6��E�A�h���^wQؕL��=�٠3�`��<��~Ά^*����F�,ؠ�{(*�_S�����q�#��(Q�W�D��~v�����Ry#@�������X��m�r��M�Cx�*`q�x"�Y��];k�vC�����4�q}Zˊc����e�E��a5�I�RX�Xbj�"^�Ԭ=���X�
��醷4�Cj �W���?.�rX��o�v#�o쩦�(y\MN�����x�(�ny�?�8J*��9y/���6��bZ��ur�cW�g����vz�4CZ�Z���85}���c�����"�ܙ���L�#����1�I�X�,��Wl������=}���H�A^nw�U����OX{��w`�j��&�K�����j��i�01ƈs&p�oczm�ܹV2y�/��):Ƹ�%.�t[l�2lROs��XRg}�8مI���؆ޠ�0��w{�*�X_� ��-�I�Q���P�����j��μ2<c�=R�]��նB�k�z�h4���v����`K�/�K��u�Ե�ya��������������0 kI����7+��F�bQF�vX��|�4Gu����q5k�U�dk?��f�͎� �my����p^��a޾����ft�ݢ����s�f���c��ż8�_M���8���]�j�T9���$�#`T�į��h�����c�����!X���V��
܉nX��P��m6��
&x��X{1Pe)�1t�	�;�BO-�Nlo�2E:�I��j�P9|�KӲv��PGp�k�ud~���
r~ ׷�}���\d�B��] 6Z͛�����d�Z��d��n00S ��}0 c����R�A��%B������$����K���Q�a������FN3Q�?�D�3Xb� ��cEe?_ʬb12/�6tGmw�Ay����/v�IÝ;�=��l���$
�U��r=�{U
�y�o<�B5e�yQͫwZ�pѰTk���h�$���b��E�F	5�-p��	��l�C���>��mwy5{�~u����5Y�������т�_��� �S.�6k@1��>Mۥ�VM���ȑ��{L�����u5���X��F{_�g���8tFs�}p�І{K�ZqV�/�0��ׅ�&ė�`�/@�)qY���y�$�'6W︰7��a]�.9�_,b$�󍅇�C����0o�"d���<,}�:a���;zOH��������(ێ�uQ�L�]I�-�j���l���.M�Ђ���1I����YL�,k9nH�od-1�+�,�)?P�:qR����� �I!�.t&,o�bUٴ����.��Z�9GF�i��Xx���
�ˏ�Ȣ���^ʍ;�#�b3�w��
�M���=�Z���YTו�L1�D���R��ߥ�"�gi���n�.��k��.!��#}տfS��{n�v���zي%�!L���1s�e��� 2��I�0�8=��%7���:�y�*G��g��+�,���
���n�כXF��Zza.�� ��J4���ۋF������}�]{�g'@��cX�x�e;ЮF0D���4e���Lb��}���A%�>�vy��v�"�O�ӟݖ%P�U�̘ٶBY@SGL-�"���k���e����.��s��^MGx��j|�H.t[T�^d�aB��s�'��59FEG�ʀ\���3^IC��\䡢�k�S���<;2��y��N>�����s��ҽ2x�\�H R!o����w�㨭�X``�Ӛl<�'�Q㴱Q}`���>���T�jʳ6+��K6��V�Khg��f��	*��Y)��-���2TA�S�wE�t�K�Oa�+R|۵�@�s��Qs'�׵	0�W�,��A6%���f�?��+Gli�$ փ�;������w����/�;���$�]�z��6�U8�&9��~C�e1�23H]������+C�x(��T�@���b�&�Dd\( ��#�H޿Kz���:���v�L)iM�N��؍�A-��
���=�۟���*�;s 4�_]<nA���vB�����������,'b�V3�J0SGz ��C��d��S���z� ��v�����,����k���x�Qgk#������Z��� ��Q�2���<��?���WC�g����#8�3%��ۇm�y�C��tIDշ�����)"�Jy����:P:�ק��[O��~�9A�5�3�s^�!D�����il�Z�c~忴��bfP�.���O��)�Y�zV�z���ӳ��#d.d��#�@��*z�|ktch���69m�c�:���M�HK�Y�ʑ�+���6��6�	��l�2��ۆ��"=ï:e�I�ϭ�)4 �w�I�q���%Tb(z�B?��윂P���m�yb�2�1�ϏD�l��*�X�ŭi*�ƫ�/�Ř?C�ư;'�_��mt�s�w�8(U.�"�����ȿ_��Q����(�hf��~V�j۽4���#��h������tT�yp�M�qR:��o�K8pܪQ��:(a�����&G�[m�_�~����[��/(�� ؝�����^��7�ߔe��$[�p��v�d3Q�\�7޹9P�K�(�O8��E�&he�͕dLv^l�F��ǌ[��7�B���*�l�,��y?�l��`��N4�����[
����
�ȄH�?f4����3�(h����g��I	f8����gp��1�����d?J1>{�
!$	�r��Y�O~T��n}���t�cy�/��Tw�4z�q��$��	 ̜�@���t��jj�'�9	��-_e��RS�cEb}!FE<�Z�O3:���m��X� Gؚ�9͉C�zh���g�A�	���|k}��CaF,����Q;�1:,��[_v�i��g�p`Ȇ�Ya�4�27�DI�-� ��Wb#��i�U^��fQ	�N�٥lm��k����K!����@�wk$�쎷2�q�|<���[M������i����D�����\M,~7���}���,d�nd>��K/#;4Z�B$���^�V_+E�-x$���+�l�V��L7oS)l�JM��0�q�� G!5z9Q,��r��������`~���vo$��[{J��SY!�����ܐ�%���h[��n�r�7n����\�D&��DͰh���SKZy���� B!W���!��hm��$��Z逦^ґ|� ���,�U9jbj �3�k��H�n��x8^��kC�pɲ�4wH��5�X���	u+*KůS]�f���5�7��M����8�O��'�մ��Ճ�o��T�2Q�@N�5�J$[cPf��	^�V��(�Z-'�����1�V�{��:�CL)��-��I��7�>�P�Z.멿j��X�}�^�N�C�!��>v�	�>
��\Qб��ޑ���*��3>��uπ2Ο:�����!�"��:R�-�	�H"�yz�9��L6��$�O'�y�0s��\\�s!��{���X�������}�$���O=
�8̐����A�1���e���'O��6w۹�,?K7��&GЇr����#��L������ �D�TS��_b��Xƕ�'Zj簺���?P$fw���Z��&�lܤ�ui�t��^����E��<�v���F��N�����K�w�2��r?��#����#Gw���k����0�M+4(�y�~�Z��n���vJX�2�J�@�57��6�|��	��2���W,݃%)��a:�O�Dp�S�,�'�M-�dI?m�X�$r	jq��̫́�Jbb@X6a�g�q��g�"c��Zx��)%��qx�+9Sk����<Pr�.N+���e=9�S���
�Cz���6�-g�I��������0o�OZ'*�`t	��^��ʇ��G��eŤ��
M�!�	l�F��R�+�8ɤ��.~f�64�J�f�����=N&�9�f��x���y:�vL~Gs�]�rbf�sTH`��� >147�0�0+�Hy�����w�a��l4P�[5M�m	�q0,o{��g�=X_56���#+����C�����X�)z���>���Ğ�{�഍FӡjE�@�r�C�]m���jS9��ڳb�ێ�$�0�K�{����Y��G�7��>)�Ǖ� A����#9�D�3�O�@��s�@{�A:�����y��2�k=uz\Se��KP�G_�oO�p#�1�67��YPmuk�|���	�bS��R�T7w�j�}���IMg�'PǱ!{����$�.aaEx�#x���8�Z�{����/�/�i뼙	*2���
CT���7��9a�	BE̔�ן�N/�H��N��['�9��L���d	U�Q.��1��4e:2�����x��~�mT�י�����N�����R#8{}�
����x�T�̿�B4�^�<:�g�°��$I������
���k��^;uu��*<R=�������χ�d��!0K�S��'��D��#�@�|� @�Dv��A�C/�D����EMΔ��<Q� s���R�����%G��S� �J��IXsaޥ6��,�'縭�v!�nӄ���T��y��p���eYRgJ����}}5�/�l�.��s�W�ϖ� �;�����D<g�,0���C�'=����`�ܽ�@H�0~k�:-!�_	r��	�)^s``   ��S��GkFǸW�E:�Ek����b��B�n��:@{���eG�*΋`g�8��ƮE4yX���)"4���ZI��W�j�F���3?�du!4m�S'������rш#���25�}1;�
j�{�
�>�?t����Dc@�Ȏ�pyض��� .�*lK9y-tE�z���b����b\�l������ջX�"�Jn��5eN�ێ��_����p/�1�np<6�i�i^s$gXZ/l!�?��,��ڮ#D&^�:��r��[�m`y�w�:<y��#5�'_0ĸ,Y1���s�B�,�0T��45�����g!�+|����ʟ����4���<�rNdZ:>�zH~ǖ��o@�6ݰ!�n$��a͹��)�i����,���6�j�����ݻA�-���\_:�A'[����X"}�F���mE�mq��z-�����ߜ��F��Z�M��IB��AQB��D�=��~ ��
�<�a-�nL3R=J_e>z��H^�P����f^HP%](�-"6Ӈ���w,�hjb��݃���G�4Wv���R?�h��D�w��#+��_`vL��a0�A@v�-�Sќ��>�)�����U��$5l��yU8�=��yP���aSwA��4��	;�/�2q�"G��e�ڶ�6�3�_���ſ2�A��Ʌa'������7=Pjl��0���bkP��}�hʄ��^�[e�}t�$`0� ��@ ����\�t�������t����։B~���a41��ty, 3=~߁O���6N�q��Ǽ%�,MO��5�cb���G3�BH��)���bq�}\�u����1�LST#�Cw�UZ+�����i��Ja���XN�`<\�3�0h?+�C������H�Qs�(}�B��h��
'�r��Q�4[�2qx��R.�1��*���ƶU��z��~Xo[�p;�}'ؗ�n�&��L���$'	/�۬c9OFz��4�jVQ����;/�#�U �%kհ�ǉ��=���_v[�S�Xo3����@���-�ޛ�v��~�j���jh]7���2
`����@�q���o��e&r/���^4l혽�����#0h�����iF? ?C��e�A��C	���6�.F u�tͅ��,\����n��rJu�y��V��0��b�F e�{�}��3�u9,�C�Ϣ�I���4(1��#���  B�f�-�6LxA�_&�5�y��;곬�zY��!H��#�o��F��h>���zz���yG�qM�b *�[�k��k6+tM=Q}�~D1��ω8��I�J}��6bd��3�@@\!l��-k���(�/Öh�B^�Z}_�cplB2��]�������O~����{���c )�ŧ�)��\�����
&z{D�n~����rc��[�����y{;}eg�ڪ�1n�~D�9�yK�����A�|�3ΥG�^�b���{e��
�
Ƭb\��07nȎsi�;��Y���l�%��#�	��:��u����.hJ��-ɋrT'+���AĘ3]R�����w�6�e|��Q�9�*�z�����y�� �}����v�`���#;Մ�(vfb�p��ޡ�{y~�r���C�����G'��j{���� �Ճ�����2��η�L�=Bs^��8��=��e��@ۭ�7s�����	��l����������i�K>�X-2����uFbQG�Q���g``.�k�����ʨĪO0M3
��FTg?no��bMh�m�#o�	��8��� ���_�Dr��x�������Κ���n��'zzіhG�"���W�j3Rڲ�
�ԠtGR/%Ҟ�����%�^d<y������<�t�p��&�.�}���:�ˉ��>�ŎS���%K�@s�՛5kK�b��#m�z����{'c>�<�y�Cc��k�1���LI�� Ѕ����'0����&T+ChR��^��@��ǹԍaP�tD;����̞��k��Ц��״"N������N�����96�����y�e&im��X:�e��Lzk�g��p���kd2һ�<�;�I�u�n�m�!%��=x���R�lVݼ3Ï��~s�$VFN%�'
K���OE/X�N��߹��/�PlG�ooɚ/-tt*B������C
�1�Α���4��{U�qG�@<���%H�8L�� ��c����Ӈ�2��vE��*0�3�͌��f!~>��ܽ馒E� lŘ��L���Q,�DV�8��*m�V;qm�g�' �9
�����L�LJ\�nf��$��X�i���3p�����8͇��w�k3U�
�� ���@X=[+�MN����45:�ߵJi��yT���w��x�(%���3��@���j�߈���5^����|y�6%=���" +�H�,�<F_C`-�K;r�$%��J"�UI�s4��|^�,��.	��FW�׵�!n	b��6WM�N��a�~�ZJ{fj�_�1%���>(�1&��JL���si_��`���B$�O��"� �ʕ�H��p�+dF�+_��`m�$-�%N�Fұb���̐�+0\E9+��~�'7��o�n��S�jk����_�z��7���h�Ĭ�F��-�τ������cEU�-^%U��%>�@z�K��/�\S?U��_�,�4"�â�jѠ�^&��T\�܈:
����%��뿏7@�2Vn��M��d��K�Jфl\o����K���Re!.�+�a"�mi/�ʤo\��Н,�n�VI��7c�҉w��$c�U	�%�>��@�Gjߗ��޵�|����4� ��v�N�I���W9Q�B�>^�"ev�G����u�b3ys��48zL�Շ���I|���)��`n��2dϪA�޸��߳�7@�� ���QN���ݔ�h�Fzyc<�,s�rlW�/fI�' �
f������h�N B�� ��+��X�s��[9��d��^�.FЀ�=�����-�s�y�����V�)?_�$e	v2%��N&)#]�"a[����9�.9;2��G��5�M�Ӡ���\g4ޮ�͎T���j��\����F��[ ��]A�T`�I$�,�5m�W���c��=��w�0�� �Aði3��C��m�u��a�,ܮQ �K��˂]��S�8�m�= �]#gq��~2�5��w�ف��5A�t5&3G��v�\��9�ݙ����(Է��3'�B�������gg���NN����|ܢ#D۾�}����ș�"���C`S���5<è�����\o���SNဇ9>�g�.���߄���D$.�ܱ����|9~��CoU(?p�!�������f���$V����{��a�?����`�Ka=�؅���1_y�U�� ����y���j#و˚w�;���y#�(x��0��ڑ���+wu/|B�u?&SX(����8W��5M;�ؐ::�z@_2ܓ��%�	Q�SI�8��M�=	4Z��_��r+�iv9���sv���#�K�D]䖣�Kg�"s�*P���K�Q��5��(��G����M�OA�#J'�jIHT���E�,���s�$,x���yR���W���jo��d�,h	.d�����~����gJno��Y��WL�8�GR��/8a�	'#���/c��mݒ}<<;�����&��3�|ѭL��F͢�;%s���T鄏��Me�Z�;��K3�ZZ����R��S�DxP���� �x�t�%��*��J��G�Yk�IK`��V�i��hS�kX������S��o����w�����i��-o��n��ڀ5~VB�	��3��_��4�U�[��@z�	#;���Wi��_C���Y�M�����_y�4�&e��1�k˦�<DQL�4O���K�� �s�U�ـj���P���^:.�$����[P�� ���:��1پ�Z�F�w���Z�X<�M�e&
&�&�25�j�ܺ��QK[v���n��vd��	� uS|��7HP��H,QB�i�vgz��<ŝ��D�w؉�i�*�\��@v��;�5��VPp	��b0[�����?T.k�+5I�5�w�ѿ�y�՞�����u.�}�+�8���5�V�h�W�{�����P�D�O�D��Wqt�>�+�K��/�)�����7(�W&> O-�}9D�bz)�'�_�
b��&",�S\����fFh�SM�&�5(n_8Q0�n�x��T��{d�ǻ"C$��(\``r-�WQjq��z�2(J��;�q�b�Zl�2�/^񻝅�<��B!�B��g�@D�1�%�m覲R��Z�;>�s���[�{{�Р��`������D�߆�3�C/�X�{&�Q�DXOm�_W�9�Q�S�)/Ud`���('u�d�	#��Z�^[۳.��X ��%�"��Aׅ�1E%��S�������f�(*��q�;+(m��=��|f������W��z�)�LÀ��$��YƊ�����`�f���f:�����z�'=Ue0�:1����'O�>96����m:�ǌ����w���"�`<D:G"#���%�3	E���������^o�O������ؕ��0Ը!��"��y�v�Z�;��%���T�� e�p�nM#+�tI�q��{��}b��qkZ�4�y���ڕy#�Օ�D}ي��?�[e����Hcg��B�v��76)�1PIӈ�1�
kB��x�5��5�Kr*���^�57��|�UKzr���U�qRm���ՠs)�U��}e*�������$5E�v�M-C�M�G3����:l�c@ �#�G����"�rW9��w�^���ET�RE4w�".'M���*Љ �p��o�5�i����b��}�B~�P6���{_�^�9�R�8r
]R�v�`�e}lO]�棛�Z%���0�~�N����ur�-�6@_�	U�?!�50ܠǷ;B����lw�Z���}�R#h�˸+Uo����m5�z��Uv��*.A��#���U�9̩Y{��i��M� �e��q�#O���*�&������9-&���:�8�Fơ�tH �G2W�źςu�T�r�U�%�zs���>n�����`�Ub�����Mr��3�K�Պc�>Xe?��9�;��
F���?+xvV��"�p@E\���R�2~�"���:j�og,Ӿ �#j�vR��U�X�=�B���bt��^O0
�;��H�H���-/��.a`���Z�^ZW�I���
H�2�1I�T�}�(�����O��g���3X�^��Z�������̲��ʡv󠣀h��m��&��+>L���7@(yv��Xj'm�8�[��۾���3��h�ʌ���M��?�!�Y6o}V�|�P©h
��}m�0�gL��^B,�E��x�����h��;�s0��`���Fo�">b}WuZ.?��3���+�@	*F)g�>3fo�鎉Iq*`�<T:��M�����
��QJPWTQ��:���]��]�Ȕ��A{���#A��B"�@�p4�'�7�9g:I2�.L�}��m"X�UP����"����
�W�!�;nLA^��]�����gQҀ=���~���E���fET�5�x� ��m4\,��])d��6���O�H�Y�B��pZ�ݷ8�4�����\��,��!0X�PY*�ŠQI]J"�	Rso��,��z3p9�v�BE�J[�-�KeZ�R���)r�쓟��|�޴���t#ᨃ�~Źs��)Yx��Җ���c�0b��f��p
v���C��Ѝ"�Vk�*��E�g+�!73ʂ��uF�*�E��T��'��))��� |���0�ǆ6���)��[w�����lt&�pk��2rV�$;���݁ ���A�_�?|���>(� �@���&]v��E�S]�W�|���|�W9';`�It��H���zb��ȅ3�B�/Kn<�F��ﶦ*���:=�n6�6ʊ��C������[�"�3g.��;������̫�\�`7���1�+�e�����W�R���ƽ�@���J�����G-���YPEv�*ͮ���]�!��6�P��r{���u�{�>F�ΙT�M�Ӿp.����>깪�e�����:��bk�f?"��Xa��3��:�����*�6h���9nS�����	�������|�
�jPa5�=S1�W�K�[����[)�f�� ��f~Ak��MHd&�Z���q�Oz�-��U4eL��1|mO<g��,[�Y�������������_~��u�����#��Z`\D��1���Z�m�Bl�}�X��浯�e��T��;)�h�w�ta��rÒNw�9y*j�%�P�(�{&��_���\�)�#�B[H�67��:2E[3i�E|�(G��V/�����r��w
�U���8=�8a2�so��d-���#��d���Xn�y`]�0퉩��.?�#I�;z.����
��'���rMH� �"��2�!Ƀ=���*Oܫ�Eu�5�a�Du��XHB:��M��yJ�m�0�5
q�; �� y-�Z���`
�Ǆ���oIaX6!�f}�PA� ����o���y@�&�c_JD1�&��"ocշV`i��d�M%�q]��S �(�����3i�����b���W@C��4);V�亜 `��dI�߇#��~3�iU�ZM)�.
��M~����y����3E�-А�&*Z��3ӽ��	p��Z���K溑��"O�9W�-� �w�cErpNt��56VU�=��N	���䉢S܃:pԯ	�*Ǘ�;�dk����
/c[G���
f����s�U<�i"i��R���U���O"U��Be�.n����J�!y���2r�S�c�";C%Њ~��������W�-��m�4��ڰ�� ���cM����2�ϼ��F}�[����%�Q�G��	A��ijn�
���&�2�LS�UEʐ{b�����iNsA����P�Ҟ'�#���%��Cݱ�ޠ�uxVֱ0_�������V����8��}P��6U��U"����i���J�S�)�}�����2��jL)�m�Q����M��vu�xr�j;�X���ːQ�����������m쮾L�e�Ɨ8X�xVCq���LT�!��$��գ�y���8U�UAw���^Gt0��5��ٯ�>
�B�>_&W����N����؍PW��Zk��[ʭ0�.�����Y���H.���*���xmO0+,H�����V��lNZ�����7VWPjh���TwH��{�x��=t�'�x&$����p��y-�I�Ҹ?�zL�	��ͣ/7
!tt��{j@G�8����G�ێ�@���ֵ���X(~�K9�Q�@�`b��Y��⤅F!�#�;�	dY�cS8���ٓ�F�	�G����Q�u(⥩�8�A�4�X�)DRԷ�a�}C`�d������Ƃ�WH �.�JV8k���Ҫ@c��-q5�N�m�
Im0�D(��j�Q
�������Ö[�3L��M��ϵe*���PL���WW������:�C#UK�q)�ax�KOYQӕ��E��OƧޕԋ ���:{_Cu���Pa>��I�OR͵�_Ǔ�e�},��A	��WZ�y�����JW���pʯӱ'�3�ԧ�"���
�I�L�����e�L�u�8��[6j�F�z`�n�$fq����%��~�Ci�`L�Z�
rd˷�n�������n�"�;>��M�վ$m��W�^��J�(j�z�Ө�4�~��vC?��`�Ɠ������̩�.V�lw��Q����Y~�P��	�����-�o]����|��jK�=��"MX>YE��;����}����m�8@�v��s'k ���(�y{�[�vkF��$s�9�*����R��'����A�ž�ݖ Ox�{��",�f�	�8J����(S�pbX����7i���{X�SPx�8ܻL^mWI}�Օy�S�/��\O%��w!Pb�3�(s�4a���7.��{OC���ꂵ�.4~넋��eK\1��V�����T�-�&�0��C֧��΄u�У���S�B�pL�Y�E�c��L��+2����~��!u@��o2��	�	f����(V�/�
�Zzǣ�P:)S�H1��k`2{�t�kl�6�i�XD0K4�b5r���ȏ�
~sI{�7���u�v5@?�. Ww1IҘ��@p�}�Y�d�`a����W}<oTT��X�2)�*��#���6������lz�3�ۆ��n��E
�a��5������!΂9cWC?1;�{�������A�u
�U$]	(冠��^_j�����Z}9!��܄�q���N�������K3��S��z܊���(�
KM�C\����7c�$1��/�XO,���P���j��
3]�p��FJ�J i-2�.>$AV6Y�%`����C�����79�jj�n��et�H��j /���������A�}�2:l�����:>��V�oC��a��}F㗍�������X���OA)���P2�)K6֨g�}@��rh�/�������/�B������ �֍K^O�=�� �J?cO��[�˝6k:�y��ѵ��Y�ÌH�a��U�q>xL��oFG�)^=N<�{
����=�	a�Ͷ��z@��K�(�m���nUU��8�(}��H�IL�]���>^�^l'�p��ja���LcB�J7Y���x���vc*�cD�)2�s�����\��#7���=Y���X����єJk{�EE^�yTޝv����e�X9vOn��o#�#�����&�6ߵ(My[�O팎�,/�d��.tt7=�K�[x^gc!���(�kp�,%˶����/�e��4\&�ZՖ���5��(7
�^��I���T�(��|�U��)�!ŝ�f.�؎�d)Lbl�˥��]�z��.�����iŋ�H��z��j=$t����G�şD��|�S#��ffȑ�I_X�J�.�4$6�4�dj*������tG��*�]2ƪI�͍P>?I��@�� X�s���L�]f�������Z�x�92���Ƨ�!1|EV��kn_�;h&�I.E����u���+��xv���:��owD$fCFY<)��m�d2fƙ��h��4IR<�Iݘp���&���*Ωl������.ԫ�S�����\��s%?�Ⱦ�n'G8ꏒ���^"b���|�O<Ԓa�I�6ُh���(	#��W��� ):��7���O3�g*�C�WJ�.��*�rv5d�F7o�Z�D	� h��7�S�ƅ7+q�3<g�mB��n�Am�aq_f��$D���&q��'5*��υ�ZE������K��MP]�F�%��kҐढ़d0�2�;V3�����b��d6�=^�=V��_[�3��ÿ��Sh&ߩ��c���90�Iܰ)��<��:�'���\HMq~-���_[V^���+r�5���`�
\_��i���~�K�=�%��u�ی�H��zC!:��kN*��� �5w��h��[�6>������K��%��)E+~�Ն�Ѻ�6:�t��Q�t?T�Jl;u�vn�f�1'�Gz�����A`c�JV$�N�F�#��_2�t��ג58_�N����e�U���,	� �}D�f�ƾ�d������]j�
�_k��@1j¹/e�.xcE���~H0�n���1��+\�}[��,�H@��8I݋��	P���k��M��j���{��۽x�B�>9��ȤI�b�V:���H*�-��}�,��G��W2G����6�T�0H�k��7S���bR�l}���"����6�y�\g������rb���}�g�4Δʊ C1�|����v�9&J�	R��k�y���.�veEO���@��P�￿�j�k$m���!{�T&�i,������5a&
�.�04����ږ���WW^_�.D[O���3�%?B;ls�|�tȕ�J�K�����Ӄ[ ˃.������`x�v���/ȩ�~]agC2�ڷ�,�	�k���V�Т��A�EdQ�ϙ��AUP��^��'8������ N!ӹ�ѱe�N*����<x9��h�4��*�t@�|
�����������s�T�K��!�*|ځ��Z�fZQg��$&��eM罇�>93�lx׋�h���5��!��|�6@;D.�Kg:&�i�XD��x��A��Ӽƀ����H����Y�N�riX��T�2|���K2�&��+ �J�@�����,�n�����D��Z�IN�[�=jV�N�/Geu��������}Ef��,�?8�,�a��I��u�M�A=��qOg��1��r��(���:~h�1�y���V�gה��>���������_�����[e�?�)	3 ُc�P	��?eH��6��ًX�z��AK���YQ��n7�hX�ժ����2����r3'��[�b���6�&>�% ��@i�#n4���?�3T�9&t�}����=	P�],��d��[EK22U�#�a�X���{�u_�74a�n	gP����!���%;��v�v��zЅ�5
]���1����xk<���!6n�5hT]��45y�TU�\e�?~ܻ��6�y���y02�&�BI$�Ҵz��l�������N�7�:��Z�\��Rt�o�\�"rcȺ���t�����5��� ���0{�P~�a�-n��,�bZѿ;F@����έ��E=���6<Y�'6�ۧ	��\^V	zaB]~|�R�&KR�6X���ƞ��L�i�6^J	�`��t�<'B�9 ���+�4��*��Q�t!,�x��3�/$І�#�Tأj�-'/�`#j���*��M�A��*���E������]1@*{uɅS�e9�Qb��$��vA���l/$�ĦΌu����v�����fHkh�-�� TWOP̷n|,g��Ψ.�v���M��`�����R͒Q!0�m�|�f�O64�j`����D'��]UE���C� }n����P�Js	:?���┦�p�Ï{�o�O;e�m��(���x�y��A$�ς^~����W���ʽ��v^%i|�[
OJQ�ٜy�IT2h�N��,�s��y �w�_;.b���h\/���CE��tQ���\�rg��(��5r0L�*��P��J3�y��߭�i���'T�k~Q�.	fz��-�Kz�cߕw8�@a��n��s�~�ۨ������ZO剪"��W'���3��o�Ƙ��߆�u�� BC��6ZqUZ��TU�{��X�?�	���)O���"�*�/wv��90�K���	���WN��B��_��P����c�]�~M�P��uˮ�W��V�-skG}G>n:ԥq��k�߈3E a����1jT=*�t��%{���@��e»��R[�$��S�M���vN^90�W�e.�dU��IN,z'<��X`]%� �Z��4ӄ�.G����K���������p�".�+�8s������Eي�@�ǯV����)!鐽��Ew�b"o�),v�#�p���y�vX�!�� ����~&�s��9(]Нe�ȸv�UޠJ���P=�%��Ύ+�x�>gHe���Ц��|�na��r�I��� ��ډ^�W*.��Ǹ�b���o��0���m��;n)l%�QP��-*�(@��}@2�~����_�u�F��q�Vyy�G�'D����6m
 $��v����m������x���&��AVe��V�L��myO�
M�&�ߕ�B���{*m�<:E��N����*�f�����þ\G��3�*�k#��o�=�w�٨��7d[/A����՜t�D7���^hwX�'��p���������ϔ�4�a�!!m�=�;���R�'����L�U�!��1�|i�X�	+u��k�Z���f�nE��\�[n���d�:9P�LӪY�c)��B�h��g�Cy!��.w�d�1&�2��j�������ΊÕ��vӍR%�Ħ�[���U�ހ-����a��O��6��M�R�j��(+��W�pc�X�����,�Z ~��+�n��/uh�.B�OE{�4�:E7^}M�B�O�����b��ѲI�)B��6y��ի9�K�/@�����5��+���N&̏ó��[�\�H���n���R �
n���c�9Z�j"�n+��܉�'\Q��ڿ���0Nm

*9)�J���J
�����������f�2V���zF��M�����$���'<}c�S!������q'G�Y���޺����:P��p�%��[����(]�����1Xab6_'�T�UI�q� ��,�� 0)��i���`f,�LQPf��6�}@fb�~v�{i�r/��'�����~��(�+�~c�&�W��ݱ������0����;@�l��2����Ę{�m��`3���|\Xi����ĸE�9�f�7�I��f�
�v��M3)
:m2�6G��̲u���_�V��QĨ�-�bLƾ,���@�"��-�h"@ɒ��/��Y^.�ؿr5�d��<��������u0*������5�Ei*bT���/cC3^C�L�j�sP��VDY�Ё5�h���f*�h��4������2!T�9Z�^��mL�/�{�7&m��}Bda ?�
7�S��鸌��mS�-���z6�!�gC��.��Ҹ�&FK�/���a_��Vd��2.@&5O�~�k򐪻��χEE#^=B�ڬɷ=��vA��O��]�����e���XB��0�9��rv�)�(5���}�;�u�}�M4R玸��� ��$MBY���3��ip}��6Lɨ �/^�& ����g�k����遲���*7`��<Ⱦ�3�֥5�a�C��'��p�<�qeP�R�}N�����ԧ����"�*9oY��+E���#���$����"@=�4?[���{?� �!>���ɺ���|�D?-�(~�e��Q/�Ib�L�e���ȋ�L��Yb���fG�x��&%ѣ
s¦.��P���Q�v^&5��7Ə�6���F~\��i�='�'Ĕ��A;��5�^e��� u��F��Hn�����*p��BӅ���ʏ�X0h�������f����`n������&nB�ei"��� �D�(ᘬ��^�Y)K���9i6�A�k25�.��>�0�H�#��țyC��Y��Nz3�%��Q��;�~���綬�-8�:`1�;�x m�V���La�D8���R��d~	 5��J�r���[��8^��r�O�MRzj>�� �]�t7��8�� ��1��$��J��vKp���1MI����=�CF\�&�����P�$�_�QT��=���CQ�)�|��j���.�)�R~s/��(��c@�����tN?������d�
���&$��<�ur�/�Y�aո��}�|&.J�����J+��F��LÉy�CQ3L�V*>�nI�s���zN�(��
O�pM�)l/��߮y��Oź�N�]��!~��v��c�+�t���~߹��!iG��RH|�\ �:4W@��MbIc�`Q�8n� qZ�t�)��,�ڠ��]�G*�D�3ef��犣 ^���ٍ���4��{�h�5��S�p��8��\����/��A��l΋�a%�}	h�X��H��!f˭J25G���l+��$���������
���8�$�	j�o���͠Q�I�r��:��Bc�|��' �vo��'��M�Td�$��[�2X�j@�.�L�E1�K�o[�6�0�jI�J���>���������ʾ�!3���ze��V�#��#�"~P�_4f;߃5�ݧ�Q�}N7�ҝ�����F"�'�x���W��O�h!��D�[�^Q�W��;�fJ5C��W��i$2$���\4�gm4(�y��Ԁ�}��?ˆ�1��ėp�%����j�G�l
@�#��O�^��LlW�e�J� �Y� NK�2򪿙so�a�%��]��&����<e,1��o�#�>�j9�׀��n��ix�Ee�D�_�Gh�-�+7����.|���ɷr�I�������<���#B&پyϞ��{=���h�:E%��Dܣv%�.��e҈�4��b��U����R��_�*P���A���+��*�� �V�Q�}���g#,���4��� e�K/�qN���o��a@/!�yP���O��D��S���g=ly��8*N� >�m��->ގB1����>��կSa�xx��D��D*�3��N�T����t7�᫛����z)F�y�G��Lu�b\�
�_��0$ޏ���o_����֚b�n���csғ��(]���%����a�^�_ZrIK�V4�gA�	n��I�-���I�Ҥ�ˍM)G�-C��4S	�Qb��D���0�%����_G���,M����W �*���w4d._�	n��W�.�9�K�z�!�$Qэ(����Q,�=<������Y�앍��
���]�>ݽKy��-�]Y�3��g]N�h�o[mvX���C�ɉf�X	:���{ey��-LQ+�sٰ�Gƙx.u!�YA[��8�	+��']�� �@����GMjJ�ZlN��K���0RԼd}�8�G_=%�wF#4J<��!���B��o�ק��9�(l���=�h�1���!��LRa�ԯ#�[�q��0m���:����7��[eF��;y��̅�[qJP��(���ǎМn�&tx�-w���\j�\i��)F|�v7k���k��cl�`���tMݒ`Q��>Px��⦑䯘��*g�g�s��/[�ekC�ȊV�G�8����P"dK��a����;(}ֹD����ǹbb�.7�6��Ň��ۼGDP<��!���g���s�%�P�"�b⧴*�.2�v".H��Vl�b��s�UT�}��~<|��*�X�20�VouaXK�\^���dPL��@�r��K'�mT�|�QG��o_��i�@ K�m 
(?����F������V:�u�7�t=a�A/�B�vX�Xl'��ݏV���:Θz��t���-?p��х�����h�%ĦF/�p��G}�� dN0��}`�#5�^���%��p �D��GD�}9�����$c��N_<��Q����UJ��k|�M���a�t��3�$��u���rN��gJ�	�ˌC\���[��e�"t���!��w��*�Z痱ʐNc�w��t���B�S�����n���ZƵ�q���gq���,�?�Cvmn��nO��#�v	,�n�f#��-�W:R����p �ݲ�FOde�C ���#8o���r��� ��jR{�ڈ�z����	�)B�F���AALj=��I����&|�V3Y��� �Jv1P%�N]�,�
���,Ajҏ��ئ�3�^��_��Rtח���I[Jhry���{C��J|��$^�/�G>�f_��+��7�p����g�T�G'�\���w �z햹L�M�5-���gpQ@����CQ�ն��
-/�yo~~��w'*�v��哬�>��?l+�e;�b^c�R�?R�_�I/��ҭj1�`�m���3���6M2)� y-A�~�\+rp��U���3��.O[�/�gܒ����ZP�ݎ��b��V�CDm�PMJ;�]�)����޿������]�Z��2�VD>�i�H�[IU�n��-�g�k�uQ���w����,{�ր��o�Q^Xh~���>AZ� ���zd�3�M���..��o�eb*`�EB�������kŕ����c��/��ه��q�`��-U��O$s�vAY�5U2\���\j���'�O,�ˍ�Fޡn4�c��f��E���t$��_�,2��N�;j!;�;k���M�hM�/2!'1V���!��w��F6d��n ۍ��K���ΰZ��`k�8w�j���<�2_]�*l
̠���Q~��\�{	������+;q�H��3� Q.��#
'��L.xϪwa~/�kU�.l*P�O�Y\�Ug��#|A�g:
�����N�=�{jrn:V{��]�� v�����8�'��_���aa_P�K�h>�[�7e/���<S�p�%��iR��H �0q
�Ϛ*�~�I� d�1 �sY'��T��ZD�¹V��y8�dM�׉�V-�"��#�P֠�d	�6ĵ���3�`�X��l[v�D��C'Z���ګ)ƣ����<�C_G�e�nEh��?�"�!��KF���t�=O/y���j�*W
Z��:v��ΐ�k��`!5�D�)���Ƿ�k�/��m�8��a'O�(���ߡ.?�iֶ˙��ĵ;��My��"�nd
�Q�i�v�8*F�9�Fxi#�����1��E�Q/�^�b%��rn���S�=`c�_ ;O���M��%_-�f1R�E��,.�'��`I��S�[���V8����]"� �]C)�Juk*��@^~⿙���AYX2�uz[����1��쬭Z�M�4|M���d�h6�ð�ﺞ�ʋ�|Mэ��Imh	}b���lC�)�[2rEi�k�lO���ɑ��p��I.4��ł�[B��q���f���X�㯻H�O��@��=_Y�C�(Zk�p��<���K�9F����}����;!"�)���m;<M<��㓗�q?R�G�`^�f��:���Uj�#w�J$�Q|S�m�e��8��"����l5����hd	��´�|]5���O��z'E����FdsTB�K��`u��f�P��q�Jn���y
@[��abpHǃ��� v[�V�D��Mp�@��뎛����.#F���Ó�e���x�6uI��� �OJ�Yأw&q�����dXgg{NXy�?!7�^��/<�F�4;(�����CZV� 3��((3��e�n�;��9��@�Wjb�FV��