��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\'5}�����CK���q������^Ҷ�à�5'4e��/NIWx�!� ��6Wr��7��)aadMKzF�<>��Zb���ȋK69}��Ef�����2�o���w����ϊb�b��^f��K���=ۇ4($ކ��k����2e%VE���6��'1}�@J�5�z"ՂË��z��ܶ�M�K�c_Njq��z[�*z�N&��������[N�vF���-�Q�0�	�z��OR�n�M�i|���8�ǭ����0�JB&�(�&�\�\U���G[R���Ȅs�*�i0����p91����R�ATQ�����3,�9��SkZ�R�P�&Pߐ���M$�����x�V[��\����Va���|u�qfR���Z�O^��� *��O,-l<0�h�k��H�����qkj;�{�%��*�o��9r�����@H�qd�֑"�1Ĕ�J�o�r@]]��LyS�1@=Ipi���g��(,��=�t��K�y�F���oM�C8{� ��M���>��?f��߹��o��7鰹w���On�?QF穧RN����Q���Eul}x�ֱ�q���B@������-�:��b~s�W�4��B{��d<�<
pjϺ����� o��O^wTn�fe�#�B$cVl83�Ƴ`��,]�+|�i�i&����!�
���s��eH`�)�.�tE�����p�9�5��R�Z#bp���������m�u��t�ݦ"->�G-��a�V�P�rA�����D[��:Xc8�3����D��u�d�N��>`��O�v�u�OܮA��O��_O-�r����^��1>٢-DWU��fo��������]
="o����v���T�/��w�Ԙ}���^��/(��4r	�0▞�|p�8&�;�R���aeVpf�ŕ��\���E�9sW~IءD��a�$�4���9���n�xe �a�v��WS�[߫��E�$\|,:=("�O��w��N�Ƃ)��S��E�K(��t>�Y{!@yM'���r�<�v�&�p���MWDy�M�nS�LeH7#
��g�F��ӽ�%WOٲ4l�|����6}����)Y;��{O�ok���r��AU=r|�^��߯�����j���bઇw�Zc�J�{cxl��]\K&h��G�%A�/�� ���k�g`���J�Q9y�At�zy�i�S�ٍ�rXԧ5�J�s�Z1�):1���)J�_������D�b��T�>L�t��T4Ɋ��KP���/(9)9V#j����閌n��/�G9@?�2��p���b�����:�����S�3�5ӹX3�FY��CW���N�$������qm�������1'�n�Nf��Ms���Y��R���Zun�y&��y~��PBV�u�Anm����L��9��5:A��\8F�t:�h��j��A�JeA:[��_����x`n���D�#V~Q)[����^L�a��2���k/�?�Ԁ��]���6�{�9�S޽E`�|��<��y9so��Z,��N�m���.��i��[]�=����s==�G���)̲�n�[_Bͱ�ޮ�-�j���U����,M��aW���lM>@D��a�	!���~��X!Ϗ���������Ȗ?�<�o0j�:�Rt��,UYd:дnm���j[�ܣ��6�9e$I�Yת3`�Y���+���Sx(h���W����:S�9�tH�ض���<1���Qd-1���:r��B�czJ�}Y�:�Y3j�^k_��c���������K��t�Z�J9`��1��}�Z�ūɸe�~��ʃ��KYD�2`�c�ߔ�v����o����X#y��.���E����� h���%�t� �tSM�o8#>0��sY8��#�$D��ܷ\��8]���T7v�3w�-f[\�u��u�C5��|��&m�jw��-ԿA���hI8� ��-�{��� ��i�Ô!_����ء �~���Ӕ:���SN2�W�TGC��NL�D�\]�>��ɪ9Q���#����;��p4Y�����K��Z�nm�0��&T�%�3U1�1&��}H�	x��.����q���P4���#9��n��T�lv�+�����*w��[�۲�t
�.x������{�txG�8�3ꋞ��؀�@�� ����ᔗ��Ԋe
*��A�ur[+��fOڠ���Đ�*PRU+y����Ո|��YR�?��9-��z8����S1lS+��>��.��Wh����q��x��y��L����\f	�#'��|�)����3@hJo�z�ED{^h��<�%�a�0��SS�YY���P|�\p|'0�@��e��,e ���!&��"!��$�r����ߗ_u��qH�]�+���>��}ga9p+1A�3���~�m8�i�ER8�w�2@J2�l����8�sy��J&}��X{:�E�>"-A���%TnB���qo��^9m}��<������R�#d������( 6&Ec?�j�����d�O�(�F�oj,w�||,!��l^�k�8�;��`����VP�~��nG�č�����O�Xʯ)�T��F[�y�"uDzK�r�=OY���>Zxp�I8O��ud[oim� -�92joXG����
d{��} a}D.�2cT�w=��h��1̓�8����C��ܶW"����&� U�D4�Å�T ��g�����(�e��XBD�O��r�O �n,"�s��:�./��G�y�eC�4�j�h5p��v��'�nF ���/�t��C7�v.���rH��׫8�+&>c�>�i���]&$����cp� Ij~-"W�v'^�o�\\�ֿ)~t�ۼ�驦9_�
(�v�*�	��n�[l���>ަ�oY�\��0o*�"}�@繭Z7�����\xLm�O_�pC���=�&;{��%��kN�T&�'q��P�<mcM:�A�j`+�S�/�N����v�^���s(41�iETwwl����GP��3�nϚ�O'�W�:j(on �9��r,%JBӫs�ɷ�c�:E��jp�-��Ax����� Xf�]/��dwìܯU��nl%��ݝ���ѱ�L������	��Ó�S���� af���q�����H�������E�Q�(� ��Ws��_�"�:1Κ�~�9�Kl�[i��������>dv����o�Ɛ��~T����;��w���5�*��?��Ĩ��0(U�-H��^fg�9ƛV�@8���We��3�b�b���6��������]#%;,��{6؝8R���m	@���(ᙅ*Ш�<�ў�uo��9@=}��'��bGz�H�-n�h��Á��:��:�'������#�HQ�;2X�s��S�g�E|���,!���X�L��
��%r������t]�-*;�y�D�r��tsw�9���t6��bY|0��zg�~��7�(�q "�7��%TɊ-R���������l�]?��}&>y�1�'1���~�Ap_q�R�r���4�`[�sa�w��7$^�Ԩ<��C�N�;�K�X��.�W��RRy���fK��s�C�UU�(�����cϏ��a$f���J]ik�P:�3�YV��A��Yѧ&�ǒװ.�E��wN��Z�l����FT T|��2ƕ"XS�f��0/2�Q�ج~�E��!�))�}Y�(���{M����S��m<(�x]�֑�Q�=����  s,V=K��xA�9���)���!y����E/��6W�5�H:���C�-~A;E��2�MUKf��<�6�`��$aV�,/�{z��Iq~�!��ӛ���nϔ���X�J��V�N��	�qK�l�/$��#ΊG1b�x[�/"p
ܷ�c"s\]�/�_�$�K�G����En�L��̾��t�֞]b'���X������f�����,����HKӟe����b/��������n�����Y:�&�����@$�r��A��)�d���VJ˒�Zˇ���tYP��U��Y囊�Z��l{��K\׶�qU�2�-IT}���Z�r)����W���@35\��H���<��u�]���y�a+hXk����)ĞO2�Q��ۄ��/�}<�	5�
��z�Y� �R*4�Q'�gpr�k�I�b����ð�ċ�^ ��q�?2�� wH��L���b�4�v�{����O����с��$i��7{L� VvI������Q3��R\�*tB�pQ�1�wFtb?uO2�u� ��rɃ?df���e�y$�K՟���ċ%��� *����yq�*�P��0O}BZc��)3OŬ?����L�E�����B[�6�BL#��zFC�;��F�r {��4��k�R*O{���i͛�³��Te�r�&��2�\�D�& ,�$����r�>��?�d.����L#��\l�Q&��n��p_��ڭ,ې NN>���ޣ�����Y�q?�.���N]>��o�~��}~���oz�432��"V*vcnpkлB�L=n��QBK������両�B-ט��sF~�	��E�Œ�v3}{�U6>�߾�{e��������!V�x�
�~3 Ǫ�!"�(y&����k��#`O)8=��G4t��V�L�̶�2'��	춵S�@���������RF��羊Bz�j}Ŷ��s2�|�:&������Jm�E	�:AG�%���J��%)�hP��r�`�V��2�����јީ��/�@�*�6[��'�K�}=94o���"]0"�S��=UJ�� 鈾d�U�G�jDQ)P�pS�9$r��.���m��qX���v"��)�J�N ;��$*K��� �΂�-k���zC�����.^T��۠�.���R�=�����>�30CĨ~`����ݧ��יӂ�+b'���;�-h�D#\�?���p�N�T@�'o��/��W^�E�%�!L��z�u���K�E^x߫��[�$� �5��'mf��9�a�`�W1�꨺H%�a~���Q�� �ݺ�xbz���+�'J�{��B{��Pf~���ۜvѤ�;ǥ�w���|��Ozŉq���(��_}�}�>���D`�\GœF��3��sf����^��A.'AUf�-B���K�t�9��A�}Y��&���l<���oY1ɨ0�������zL��ej
��#�L,.��J�嵰#�����V����qL�B�N��l����#�����ZJ� �~ڳ|�(���_�`v��bO��t(� ����,���W���ߠ�>N�^��(i\��՛ �7��h��W��=6a��e�~��r�ۅ��UX� �1ў[�n���b�/�D@w�+�JH�1��S1)��2��{x�I	ͪs���ڴ��V>�=�B�.�N��Dʰ�4EA����#gx;��ZR-i/g8�B�;J��v��BW����)b��5M��Ⱥ��hf�60��;E�Z�ɛ��"doj)n�h�QӎX���(>~�&-���A��-�:ɰh�
�.�\u_�j�w�$a<g�K�,T*���I���޸��+/8��:��[����&Щk�Yj�X��MKwS�qo/ȶ�������3�s��F�g�R/�G��d�L'�v�271nn��8;�<ʜ��IĢ���3�@^jl���[�0��>��R�\]��o3��^�b��ݓ9��ZHm .�.QX{�?�<�cqgs������vMX����%$+�y��¦���M����Y`aC$��\�*�w7B�l�e��N�t�7�S��*��Q���;��*��ߕ���(�T�8y飡2�ڮ��vyu�9
p���s��0݄�Sd4�p�%~]�A6 ���no{�fjj�g��Ձzc⨔�uQ�&L'_�2;���qY8�|1.;�T�9�OZa_Ba
 �C����D�d�j;��I�=;+�=��$e~.��0Q��x�f�#�	�7�����WȰ,�F�,�@N����_W�Q�ͤ�s����*?"�+/�N�*ܾ6��ݰ�Z�HwoÐ���F�.��~�	�p�2�e%8�,\���'KD�3"w)��Kj(I�Y��i^KP�Y���h�Ik�,���ӛ���eIt���]�ԫW��б-P5�:�Gi��	�N�<�<����� �4�v<A2��z���6�|�e�F�P��� ���V�w����rW�?iN�\�`��'�����#S�A�96>k�+�g� �=,8
�r���qZX�x����sV0w|Sݕ������!���y��	�-��`v�7g����1��8����$��z^�$M�xgcJز3�j�	-���+�� ��� ���-�������+m!-r��Xг��uǵ�����:Y�OS�x0���}*�E[K��I6��R�JL���|:�N��nC���~E�c���rW������6򑖋�����W��`�,�HA�J����R?�J��'
��b�����n�Q���F�M:�����K��+�ɢcRՅ m9�Q#�v�@3 ��t��m~�\��ZƱ�z����||�]�<�&T~Ev:I�HG�[�>��Y���>���@5�^%&X>;�����:��㊙��늯�tR-�UjKP�v]��]�X�89>���q֘�g"~� ��jy*�5!Ǌ��=+e��Y)�cM�{�}Gp��T˚ͳ oΕ_�.���GC��Br ?_��Ѧ�Kߗ~v��lP�LĖZ^��FVf�� qx�������9	���	�ߨcHZyȐ��˗1����r	�__���U �V_&p۹�Q��t�38l}៍�R���.����P�9�8�Ѐuڗ��p(���jQR��%�-1ݼ���6C�?�T︈ET���=���ۍ&��a�-��gH�@�=�aAւS���c&t��O�Za��m�������9"�;�������AV�M�ԙe��e�˷k�}�������۝0��#epǐ�%{�]���8�po�A�e����c��-m��!��qC���+�/����1�9k���%G����� �V%^�-�Y�Ȩ!y������q�Z*��	Z��Q>��To�k]l�bHُ�&�z@�x>�qR�(y���6mc�h�2o�ܧ��|����+Nn�A�L8P(I�=ـSv&�����uz>�f5ItH�m�5&��()�[�:�k<J,��"/}C�f�?$�N�TJ���6iaG3L�X�8�ql��UKL�Ql��dQ����~��0�-�k�L���}νǴ���
I����G}K9,�����jCD_m��[�S�N���,6r��F�Й�m=��`.C�ǥ=�����Dk�ʆ�d��Z5���k�m��H@7��h��Q8F�L�h�H� �h}���r�O��~��4��Cf����]N8��֥pP��"R�4�s{�7��<}����ʚ��Z�V�N̿p��=/DǑ�A3�]o��Xt�r��pd���9��2�h�|�_��r1��X���_�M��p�H� @��ϪЕu@�:G+�G�d�*���l�~����]�#:V��A.�V�&�,=�B�Ї"�"��m�GԦ��p}�����wB6�g\�l�GbfWf�u�S�`	Մt���siQ66`�)Q�h����QU��Nl�A�L�0h�M]Wn���6�	 ��Y��P�D;\��$4U�>���`s����
 �V�p�1�_�)waI2}�Wm��}��c�w�f0���KS���������i�|K�hU�}�f�Ȉ9�z����ja����X��!�E}�7eb�nY�!��c�C���l�	.� �U�Rnv�?��}�A�D{=륉��
�G�Sx�mEm�j���۲�j���s�*.t�ͦ(���f㭻�r��]�'t*lXa�8�H�<������v�M���Î��@oX�ep�e@/-��r�)[S�Ee��0����-�*��0Z��9�'���j�2���$�d�� �c����bŬ��2O��w�ٰK��XeK$l<�$�e;�H�?鱆8ſ>�h�t)��!���ٜ`�l@7�	$hN�(oz��'�,G��7���:���Yj�C^�Y<Hb�QU}���w��pot��] @��s�^� �ǽ�����҅���NZ����Wx=Uէ��E%怴�魇����G-�7ѝ�C�Ʃ6�2�w���Gi������߹]a��-��.�M���WY�aL]ۭ�_@������7'Ρ��>�uP4��/��j�?*�"w�U�����`~�,�����C=��om��6vA�_�oi�U�/�C*!��P_�S!�^��;��9�ls��P-a[��r+���c���`�X¯�tŎ%�s��`Y���R�R08{��D�_9����I�だv���h̍lz4����i������9�C�������,�n�-�O5�3��&=
'��x�����;��Ea��� �@˔θ�>Jh�C��1ls�H-e1^�fU��I�׉��K�%��]6l{UO�Pq�X���n����j� '�Ge�>"f�81Xj� ���֖!�ם������5p 2SW����l�v�S��ׂU�4�7�7~�oB���Lo���:���i��^��\r�B��pʎ ���:D%�D�ex��Ɏ��?���)D��ʔ�&��"B�LMMA�����s#to^�FU�CN/*�ᶑ?��:a�[\���b���J�%@@;���Ρ���:F��V��}�~兠R,6߃�%yIܽg{(����T�%`~pc��b�w����S٤���L6�e�5��S��GI��k`h%�Bg'�}v��$jeŏ��]d�_w����"�۰]dĐ-��+'�~#7�#���9^���w� �H���
W�,)o!!%���b�"v-�����T
:��E�mf��^*�D|3��6/K��ߢOϿe6�+����'51c���4�j9�i�9؀���V?:�(7���N�t3��nnT��j?$�&$Y�0�$�A�k�	]�Z-F��8AV�d����߽��֏�Z)X 0e� {.�����_Ύ�\��@7�����V_���3��E+c������03�W��Q�����2�_�C����>�O)��������c�]��%{�r�fQ���s��V��g	�p����!�/��E�k�2:�j�"R7-3j4.PtNTvb������U|W}l���^��A,�	���	��<POwU�y���Q}��ÐQ�G��5��Q����,$��up�9ڕH�Ў�Xy$���yke�?NRs��=]�.Z`;�m�	�f�"���ż^*�5Ԟ�Y$/n�
�����ۀ3o)�z�)�ehu1��5\�Uo[�<�3��B���-op�K�q�I���Ny�������:I���ޔ�wg'`@����]��CkHSsIh�ߊa�'^N;ǧښ"`��3ВT�h�F��ϟJ��i���|}�z���\�p�:(��'q	L�ԏ�,L���t'���P��L�x�y���gR��������7��r
�|�^Eh�1�h�VO�����X�N�����m�ݘ������V�
d�*�Y^*t��\�_�ES���փ%�_����A	4��p���
�N�#�����d�>T�(��*�j����a�ު��vյ�����Y����g�7"X
�eOH*���I�uKd��}�\eA���O��n�9���F����_��U�u�)��`bÀ����6L0�'.��d
�ϣ�X7���&�����'4���Y�
��nx����/"���4eYGS[��V��<a����;�85�D��"f��>�Zq��R������������3�\WI�����a	C��j_�b�*#���_�jM\��6���pk5�\+�sg����!�AG�&tGE;M�_�R=b4�90���g�3ʯ�	���Yo�pN�v�x��y�r�*�WU�n�^���w7�/�Y^�y�ȏ~���0|[M)��M���j~=�d�s�J�^��o3Y|$O־~�Lf�������)���J۽���&��Q�w��e�V�6񛟆�ǰ�kT�O�#C�ǯ6���M��9����[������="�a�����f���a�%?�Ė8ǥ]��\�}�?~�5�����Ap%�e�0�9F�P�� rA0�aD�]'Z�~n�N�j�(��/ T!�a�{F� �����o��m�2���s�����ڇ#i�'��)��GjmMM���p@��Q�w'����5�`}wH��Ε��?��(_���^�=��AX�Xc!4�3Q�5��b��Ӆ|F2���oz
&�dJ;�/D ^c�.��P����¬C|��ϙC��(3�C��q�Am^��K�g���#��X��if�s�7�Mh��\��ϫ�$�R���d�x�Z!>�CՑ�-��Ѝ���<+��M Dso�A��70����l"@�y��7�<ߧ{O���6x��=�n>L򁄞V8�Btz����"X1�A����^��@��y9�g�h<�D&m�)=�r�$CZ̏����/1+�R?�ns{@�+@�&�C���ȗ�j�wT0;ur����}�Wdvv���M�A�p�)7�� �0���Ĕ'�ņ�\1TI�� R6z�m�V:t�~wϯ���,�S�:�&�u��}�
S��;;ƹc��;��N��^<��������sh�|�@��Q�˅����<Ϝ`�S���͊�Ԫ�X�Ds�H�����С�;8��+���[:�Q
u�Ds�#5�&��~��z0#��RD|�G=|���YDYE���q�����ݼ�xv|n�σ�W���v�;����{?��� �򎆅$�6��4���!�C���S�U��"�_nY�	YYT\����}���a*�XW:^o�P�I���ӽ2��4z�eU,�X���/�ט���屟\x�ܹ���y��ض�%����k�+���d˕ �e�����d�ǄoHā�ˡ�o�`8���k�<~�"Y�Շ��E�U�Y�Y>lL���]q�q ������{���*U������!a���4E�/�j��0,� \ؓ���z��&����f�y!�WFSm����6 I�6rqy��s)/�ɠ��(�Ss�L���-��Y�ڙ0<�R�S*���}�s����,#����;	�X$\���J���d�j0���(R�"!�_��ñr��$o� �`�ꦏ"��9��Q�����.@b�10n��X�͆�Y�+��ĕ̺CXJ���m	t�GCj�׍Ϸ�'N͋\չ�x�ٰ��04�r�7���iV196�R�Y���<��μ����⪋��Kf[�}Ǡ�0ɰ��҃ôs�<�vG���u�7G���/�A�^;f�225rc��	�t�� �r�j`��}bu �h,i��|���5߹WLTT��)�����ccR��ī�(�<�Uyǒ׏LG���uFE���q�lW��s�9;,&�Fƙ�1	z��vC"���}G�����)�JMa�`4���7�)+t�z9Ku���Ɨ��ۛ{�m|X��X*��ʥT�sD'�xYF�i�\P�G�w�S	/���Ӗ�y��v�1Ny�(���@��^� ���c�ZuZ�V�=P�D�lx鬣N��H�'��&{��N�e��gꠒ��6W�G�^�#n��\Cj>�F�7�+�)-�Sn{$�Qc;g*�W�^z�5�P�������T(|,�	��ʧ2��e ��zm�l��^�
>B�qpXEǙ�g��2kc2�'>����4K��q=#�6�"f4���KY�?���L���K��ญ���,���hI�=ɴ�G�������a�њD<t�9�{�WR�ag��=��j]�8�.n����߫��5�������!�Q�-�y/��hFL6���W�8.7�/}`�_�wl�e8C������Ҹ�A�����U�v��ͥg)�5x8�f��..q�%���6{&��Z��s�D�68ЖD�@���$qi�޸!z���H�u=S}�+�뗤ˆ{�ƩŵfQ�[�\��"�~�APdYAһJX]�dE{���Z�0��i��fcMy�HgJJ|����'�ˆ$��G�l�%���n8���%eTVL��G낳�|�c^Iy|kٗ����g���AG�[2��L��z!z�A_*�b�G���Ծ͆��+��K��6l���&�ud<.ЕOo����K �rZ_���72�?���Ui��gg�`	�%婒�zo)H<�A���^�N ��ya�e�͙��!P��S�8�h{��P�_π �ۺhT�z�?PT#�e�ΉoQ}״�*���j1~�5LH�4�6]��HZ\Rb�|�����dd�}�鴪����t�M�+/����m�{4���e�(Ј+�B�I��я��T ����Mi5Rs����e0(���jr|�Z6�.g9��	�.�1�ٜu+����D�4�k� J�ള=%��tt��A��f��vҧ9���2��>~�����\���A�!�H$s�44l��ȯ@�K־��:�;E���X-E�QѠq�(������^4��(j�:�ä�7<�qaW��.�> ��|���n?���.9����Y����o���ZuX��M��q�`+<#��׮�E�p�&%�p�"*����8�誖ZD� ������h�HPP�
1�\�����]��8��Ͻ�������B��%n4ޯ�~[?Y3�BAU��G��A~�"�����n�>����
�D�V<O���HޱU�����>�ג \B�e��Q{
�g�n�żb[�z0|��1g�ygBU�����x�s�~�=8��H��^$�\���F�@H����)��aPxŋ8�����-�����#
�����v����[�<I}+F�E>ā�ߖ1̲eDI�ZU�
����0�x�,���X~I(�?]��� �<�7E<@,����cxsz�������!�'�A�9(�k6�h�"�/��󔄤�Ȭ!�n*������`[(f�1-�`O#�A!����@�ٍj�V�_2E:�z2%�\�"|q��d��l[Y��x����*�O*$�H���tL(������:��{ �f�P+*I�+�H4�d�����Z��-`��^�L�c�s�T�x:>�?�> -�Fb������􏰊ĹzZ:?+?Nj��:�۹�x�h�&�ECL+̃�@Â7��@Ix����7�`�"�XЋ���<���=hzH.�g�
�6��4��^�:��|08hq��J��fb�<#^[g�ɗ�&��� �����NY�`��4c�D|&)�=u6(ߔ!���5b����)��J�dB�������G��KEJ��c1��nt{���!�<vDB���ZS���Ss����ϙ�����S W[�擌�G�Ч����c�e����Lr �K��N�V���a05�y�$��HX��)D�a�����K�Ǿ�-\�I�Ȟ�˳�#/���Ypp-J���̿���o&y�2 ���&퀇A[��m�Գ~�[=�*!�k�93n�m�9�aX_b8o�?���p^��i���^�n��ކ���⓽ǾHgA��d�q9�|`i�BZ�"��Z�Z�0>@�j�"�GD'�V�Z���>D/�I�TG���O��*�uM�OMl����;곝�v"�Q�=yPg�$gj����\o����˧V{�c:�&�vS���F��V�L�f�� �ߡ��q��W���E�!!��ʅ��#*&���������u��DT��8�À�)�d�r=�9�oǰR��j��\D�D����Y9���Y[C�_bc˝�9�X��o���U;n �2q6�\�������1��%� ��������pq�ZQB�ʞ4�q�t�����T���Yr&C���-w���AA~s�K�ie�@�۬��3�8!E���K�RJ:�x�o��_�s��(h��p�w���W�{�(KB�\<T~Kv�9�?�ᣧ�&!�q��F �_�k �Kf���IhWZ;e��L�L�n����q�'���	fǹ��T �Y(�j�c��NŶ�I����~q�*������ܷbe졹��q��	j�;���F?#�"_v^��	��W?H��5�c^�#�Q��Cժ���a��f �&0Ǎ�+����o�������Txƹ�0>0�T;L���]�,]+���W�(󁱮�$���*��:�E�'�4v��\�tB�Օ[��Y��&�4�ӝ- JC&��v�5��S S� 7�(��>�︝��v"��럝�S;�����0�8	c�/�B�gwx��Qʳ{���]��b+�e��-�{ϨU�}i&t'�����,[z�x�P�8)�B�p!/�ǒ��L�ҁ;G��<��̛��~"��]�Ё3�w���si��eG��"�"*����fSt\�
�4�_��:?V9i��F����/e�M�5��!��-��`��؏N��;.%�� rYd���cvl��z�������<%髃�A��-_��?�����<�W�{AH}<�I�xW��Կ�E3X�Ӧ���6S Pwc��5R�c���W"ą�n��5�x+�;H�>�%��M�? �2��5 �"�x�h�B���D�ft�y�3�x�e�L�Y���TK�!����%���,)��Z*�r}F�8�bncYթ�x"T�`b�|qSu�<c��/+� ���(qz3i�(�sl�/���DR��&i� ?��z%����Ƅ(G��u���ce9y�����&����{� `��ƞ"P�Ɲ:�nȳV^AT��|�� 3�{cl��D�s��I!|�uJ-"%(R��z�#�ȗ�g�P�l8�~! 	Zvql@K6),f����}�_l��r�����'C��i�= �L�X<3%�V1��M陆a�TD��������F�ɩ���ȭ^���F�?��3�����O� �1����S*�ViZ��?�}_�8h
�H������7c�Y/
._d��ˮ�2Қ�9'�&>��%bǸ��k�.��Pn,��y�Xl  �M�u�+Yw�Ҵe] K_������H�ИE#&�������.%�c�	Z�s���OD{��9^�3%ޘzڀeY:^
����c!ɒQ�4k�:��>4<�uP�1e��(#�����~܈����A��$��y�AN���=�-��}�k�`�4�~[l��r��T&�h#UX�0��D�#���U��'�ԁ����_�=�b)����_=%�x3��'8U4t�7E�����G�|��I��3M�WE�[����{��q���Ú�/v�A�0sZ���d��7�E�����ʤ4��2�P�
��wig�j�y��}'a��La��� �op&Б�k ��i�:����A�)(J~�>K�m�~����L�(F�b�`�g*��C679�s��!ʮ��.��*А��j�<���2��D��mb�EMr�������ͧ79���3��ge��dV�T�<-\���#P�C�P�O�-��K1dH�h�*#:�+xF^�n��I���^�gk5{����z;��y�Dn'�4�k�m�:�p	r�X��k�B�PO��ꁇ��:��
Ȥ�Q�w��<|�E|3��������9֮:��85�zA��hd�gj��V$��Y<�����+�H[���P��u�'��D��aIM
�05�j�+9H6-d2����N�U֓�ݖ�1��VV������q5E�g&�6| �N��C�քS���f/?��pY���Q�w7s������o�%�Á5ɳ�)�ܢ��Te�t��&��~\'l��v��NJ�."����l]fj
�&yTv��>y�7�v�Z����(AF�@�2�zb]!��e��	�|؁vV��%7�_����Ц���FN�ƟL��A�f�ލh���8G��n���gз�Lѻu}��,v*�3�}p�M�L߱��R�>�qQrRؒZ|��%\P紕��<Ү�˄�b�U�n)\g{���@`EABZ񳑠�)�[%�WW�y����ąw�j�V|�,Y�0D�Ed��8(�3 �밷��"�YuN۬��}��®0������ Ċ���*�gL_�6�Z�� �P��{�KA�V�47�WVd����ji�c��茇93n����y�XgN�!�I��4�Z����>,z~��Z�u������JW��S�#�7�*�}1=T���8�~��03h�T�����x��ߨ��f�|]a��IY�JyDk�Z¥�ph���3�	ɝ�ץ� +T���0�Z�݃U�c���j�neZ��>�CUYt�K��i8Z59uYak���)�1�	���4����1n��rd�9o�X��i�=S8���͝�$�yODH�4�f��Q�?e[O�ۍ��S�b��8�28�l��^���0
�ugܖ�)��b��O�"�p�C�gȼ����<3[����Ɵ�;��-zW���cj�u�;��Z���
1QK�P�Ӝ�M(��h}�3��:�]}b�I&�;�`�{��Uժ([sv��@��!Q�DPa�.����,7��",.��!v6㷼v����-ȷY�*�XE���>XGF��K��>ZUe.\Զ듒�I���l��sC����/��x%��׸���\9Ð'�kR�P�%[��7r��Sx�+x��� �	P�u���o���dJ�>�!��[]���捞8.Nzk�N��ʚ�*~�����|�O&����	�m=�ŦX�2�IӘ�HSM�OY�پ+:w=��D��YYt��Nd��c��\#�K���yg)0�X-I�De		r:��K��yF��ٙ���|C��l��5g5:��%�Ǐ�j���1ce_���.��;�ǾL� ~s6������O�R̓�)#Axvh�F_���v�}
ۡ?8f#ʝ�_��e	{q��)���*��_��xj��UE��r�U������z��>��g	�Btw�1w���M��:�բ���I��j�W�{v��}�Ja�g�,e��|��S͇i!���oA�x8��uE�" t�@\�G|[.&˼����6�N�&4��Sj��C��Y0|w�H��h=[|�ura� +���	>�wN���i/Q�F\�;��^�h�Ʈ�WM�*��%~�U��$쮌��^�����e3��-����N�V�|���x�rI�a�����+�O�j�f�#��o��:���7�&�#�X����0"j6�/�y>��a�0L̓Ou��q��ׇE��h%�?ȭ�(�3�۸H7׏�<��,u&wC��>����e��Y�"�C���7��ę(�Q�����v�!��O���:�9P !�c�E�,	y˒6�| k���4'�lNh5�J?0��IכYO���.�^ϯ����g�i�oCA�~��gźt�݄��^��Kx�=���\�.C� �.}�r��X��F����Wź�`�д��ΛK�^҃j�O�hY���	CY����) ةCL�wuï�p�@	�����V��e���>0NL�e�G�h���W�4ښ��c�_�I/uR!��es�H������]�ޗ�o��|s�')��0�����=��H���V�q�  v����;��GϤ"�3�Y:#��-��v�o:y�����>"8Ff�0ِG�=S|�#b�7�8Y#}V/�nV�n������N�
�45�-�PD�k�;P*cT!v��HMr�G�\��iILD���c��K��nr�'�T)gG����"��y��&�Z4|9�_�L!��X�����xs�s��ϭ B0>o ����]��6��"������W�Zʛ��r�����^��͎
�q�b�epcP5U����j
Jޛv�i{k;S{�d�ٲ4��<pvw�%^N`�j^;n�\̰%S;��sq3�Mup�V�ɘ���jݶ=�-UR��*͢3sņGp��f�������}]^�n�	'�2�{�>i�x�\2��-��/�x�,ی�����]ƀz2�0��)�vâ�Q�o�/�㥱�{93��> �w�э_*j���[Q��v��X���*�̐<246#?���`�YFϼ��m��`mZ��^��չD�@kC�lW4��(A�M���rdv��Ò�#�w��,�l	Ak'�Ҝ9d���[~�P����^���UE���ޡ%dsr���}�[nU�#�?�X�K����d���g�����I�U'��F��B�lW��e[0���$Bp�`���a��TP�*�@;R<���h��n�b�(�����V� ����$��n�V��ܩ��AۧJ��v��^f���E(����B������zϖl�՚��E#�b���^�s���"D>f��p~o����u���oe�c�:��(m)F��
���?O;��BW�fZ�.��X�+?h]�r�L)��n���j>H��+��{�o��~~k�׆u�K��Z��.`&���nKt����=f�LW[¶{�bA�ʹ����jhu�i�͜l�`@>�ϒ��7����L���d[���`�+ǿ��+�m�<1xJ�6b n͓
y��	��a6�������ʺ��¹{Q��e#��B�DwI��Q.�6����q6T����5���y!��]
5��Zg+�J���n}��,8�����h�37W�?�x��UB�A10�s���ܣ[\�k'%n��vY�����.�BV��P��u� ���
�qeu.�#��u���j�g�Nr�(
Զ��X��εg�ْ�d&~�\+�F�v`�-	885W˝���� G����G�a����1>�1P�yr�)0s������m�.�~��J6CW/3���nwhm��kE����;h�$w<��x㪣���h��e@���c�7�u��Gm�~1(pӝ�
�b��g�:��{ć�契����"��[w
�rG�L�mM0N��ʉ9��yEu����p�KY�_��HL�- ؕe����f3B̎����譡*k}�z��<	����"��K�݄suAj���3z~8ɳ���U/�p(}o�cQ�U=/*y�{�e��Y2�'�
����� Fj!2$�C�<N�V�`�V1�������#�Ju�hs�=�ys�A���c^�4'�IS��q�/���	b/��!9X�<8%��a9Q8�n��8��������
N�������Z�wk���Ȫpt�ד�z��Ik"�V�T@2��(.�����禳��:{mE��2=	��_���jz�7��)v�+?�C��C�Db8����������+�+� ���� t���<�F�@}���l�G�m��ʑ��fQ>,ҧyq�mr���I�,,�����Ԟy�sovN̂Q�l���l.'��J�^J,ʩ��쮒�r�	��c'��)库f0'��Ĉ�YB�N��$��o�x�v3�3]�t��Mi&�@�I-�@��#�G�Hkd��p��ǿL/y�V
М��~O��\�Pʣ�B��+p��
I�X����n��N5�� ��\P�.��gVA�|�'���ݯ]��2��;� .�{�wh�[Y���j�2�SL���D8|��%���ܒTh!���ӝ�.=s���;cT��1��B�;zX2�ꮇ!���wo&/ʇc�b�ƛ�%�DfQ�� ���,Kv7_A�ȰM�����lG����y�M��/��MY��9�l"ͪݖ� �#��䏯lĳT�Jx�� r@�d}��a��	
�Z��m��B��h���0�k�	��Kb��\��I1ȶ�d��fY�U?v�BZ� C(� ��U��)\��GxxLx��νJt)B�҄\��Vɮ�^��@5�A��	��2��2���V��[�V���\k�jgǏ�Dq5�QR2iYW�7��Y�k,h;'w��tl����	&O�F�7؜�';�fGh�<�s�$�����*֗�o�Lf�v�'V��e��^��C�}+�U;�r�$��@�0�I�a$i${�z?�v	�_�X��MO��p.&U�ILG1�4O�x�(&!\���$S~��<~��-�Z��Ij�AÙ� 	�k~	�"4Gg_m=��;8�Ĭ�>�Sp����� �	e����{�@^�M���|C�I��KW��i�͌�S9U�֖k(���kq��e�#B��$~�<�f�U����R���s��wA7d���0�� (����p���5���l�p������}���9�<}��.�����
r�]������㓿�]ʹ#հZ�pU~�������1� �d+�Χ�`�Tk��gK�X�>Fߓ��'�q[��Hy�}���-�6����؅ź0n�<&�R �ϴ!�HC��{�� �1a��+�j��Ҍ������hO��v� F�?��#�0_�.�r]'���$���w�:z���~\2.�AQ7N>��(g���ؑ�����v��� ����f�ξS)w�%��-�<���}�sҪ�;�M���݂��0�P.��m�̒����b/�u
��l`/*q����#�X�ưrk��	�M�Z��ͫ|�u�(BM,@HEW���dl�� #���	@���a��(Yy~��<º����2n��������;:��M�B��`i�Rń�ԣ�m���b��35@5T�O�����=6������
���^qw�%���YAS�
�@Y.���|3����ŠPc��-��B?��(tȩ�Y,�,��ζ�	G� T4��K-�u#KNM�۲$�ϙ�/��M���JgG2���,�E��ir�d7]�ئc U:�ò�'a��c��G�L�b�7�L� Ea�k�h?0���$��4*�T�W?�t�7#5�k�?��3��_�`��1�sִU$�* ��]c��n^�0�iT�����:O�K���\��4�C����i�;�*+�6��XK�[F���9eGr�>Hv�8ZfB��QaDךl�=�*�X{��\��S�������w��A�@t{��,��p{�r�v��Z8QT�_����g�dN�*�|�(����*�"L��ZL�AQ���!.�������s�vW��@#��׶IIT�g�8a�|�P��D ��p�0��#����,�u�t���7*$� ���R�%�3�:sup@��P���8Чp��?*�0y$�4�x����g�E���k�$�]�X�X��A��3��N34~+�io�	��6!��s��-0�b���"%
7b��޷��q�K���m���fJ#�i�K��O,y�N�[*��1�̢R�עYlo���R�Jv�NAN��0qH.ۻ��
����Gd��k�<Y[C ���.dc��9��$ϛ����	�/ 2=�U��(���@\Ył�RO�R�� �H��0��̄T)i�K��wY�MI
O74�����}DU@1��5�nss�|C!��j8�]J�v�����W��`M���?p�W�1����\�������<��X��FV��;M@K�+�Ā)��D��g�&BMW[�#�J��Y�Qv�3qq�U�ªF�ۜ{�A���Q��ϐ�����]�\잦7x^r�jf��F���N0��U5>'�g�MY3q���g��jK�"�̻��D�8}��IЄRWA_"�*#�
�w�m1`J>_��*_��*!X�5
�(C�Z�;���[��&�ñ�;���y'*���}C)�ے����-��2��c�J�a���Õ���X, ��m�o�-��,"�<M˸})1����1�'��3�(y}�(gPpGΙ쐣�7!����yXH�����Ϗ�X:�J(�!H�Y
T��)��9í�έ�����������ÙT�m�J�o���F��+�����J��U�(9�H�{�����u���ŰL�!�B1��EѶ�6s纷5<�t�)�dz���6^j}RV��s���r4�HR���B�k�$���y��M��iuV!i�t-Q��g�a/��.5~���2��]��W<�[��m��Xi5~�:��5�LE�V�.�G0��O�ޤ���I��x�%Q�ڀ�����C��$�DT���I_ Qo[*qg�Aa}��Ȭ��Fdz����O��nzaL�~��\�mm�ы��D���
`���X���f���D8���凾�*4�����4���.��*I�hL�ge`uu����g0r 0q�#��`h��i�h[){����f!��i�4����"#�MG�Bg���	x�Ŀ[{��2巬��)��|�����H��Erve,=�em�!��$��7���<�@&w�$7VS�������Ӗp4<���_%KSKwh�k��