��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga��E��U�z�����
�1cv⎣�/�h���ʀ��8����EE���<��^Sc�Ѭc�ߴOG/�ۦDh��P�`����T���uz*dIE��Q{j�z�y'��<�CS��Q��=�@o����L��	���l�K��om�驱 ��葶&&�C�At��+���}�s�;u���,��<��gQ����kWa)'rQ�P���JL��lW��W��D�^��?�/�ٲn/}^?�b��<��8�ک��L!
*nԊN�nΞ���7n�`ʎ�~�{���A�l�b/C��&��`��8Q��˪�j�� �k|r0�#�ki���_��a�4�T�N�=�M�m��Ź�c-߱d�����:�3.����.oB3�;�е��QҠϔ��b��eUnP (u"CD.�����V�e����]r5RAb��[��Wnx�Bxs�w2n#�C�iPA(��hp�����W��\�:�xc�*m�ګ�`$��2�,�Q U����ԟG�ʬ�uhܞ�Q�u��G�@<����&�By8�oa!�ʟkb!��C3��'�L��:�|׷������:Q���6�c
}�����F���?�]IK����,�h�L$�d�fYG6�S���ڹ+2���ɽ��l0Q7�7q��g�{�n� ����� �w���C\)t�wOb��гӠN�����L)�C]6���=��Vѝ�b��/���l�_�A����F��郦Fc�Q��jAEϡ8�{V=o�o�Q�z�S3��w�����Z��\{�z�� ��Zw����(R������\CW�F�xv��ۀ�M��d� pȌ\Q��u|X{��3��K���2S�f������srAxz�n�v�^�����m����*}��} 9��DI�kZ�|�A�?�����_t��κ4��R��I��tN�\U�D�E>�g�w)
��ۼ"�NX�.҅N�{a��ǻ�@2�o� �͆�u�J81�}g ƣ�RE��;b ��q���H��^�g;Ԋ�zf98��KR���J[���Ȅ�kzc�Ynlo���XG8�%�; ��ݒ��(5��f{u�J�*�&���P=H���C~~K�$��썬JC�#������%��B���D���"��-GM��iW$ރ�z�����PȢT��V7�]�Y"UhS=�On�����N��w\&J"�|������c#�t�Mw�1qZT�AC��2�](�c�;��R��<k�W�'�
T�X����[:������d��
��Y�̢��~���( G9O���y����0׶YZ��\�:i� �!p���f�M���OY#�̾gT[�g��7���w���/e!��2��C3�6�*Yϐ��*�i־T��'����F'��;�~,+�L������`�{���H�@3sZ�5�z'5L������*1���������,¹j)���j�ߡ��>�D�n�u��5o(����*�PC��r��V4����JT�IL��R\'\4��_z'��k1�T����>cM�����(�N�oJ?.	��P
Pi��7lx[���߹~I�J��[HqC9�Ux6��Xa��{��=����9�!4��b_��1��tI�	ߞ3M>����]qE-qv��Z�jAe��2�Mo��|���nL�+:}X���ش�|��L��\d�b�wR�AS�gM�x<�y2���I \E������]d�2է,�#�?\��nޯ��&�g�:���,�k�X`��C;=;w�ޜ��XUUme��s�̡����5����ʥ����*�!Yȼ�E�]�S�(�=;��DA|+O�IQ48}C��fǶr���H�jT�<����K�u���7��Z���:�Q'�c&�<�R��rR�{)�w#�c	KV�_�|M涒eXL�fD?��|fH�Ē��� ��BL���tZ鞥�Im[[��(Ƴ�R�� ޼�p���'_�w�CBAƇ��'BU��dd'�Bޕ�u
;�)��̀*�p)��,�]}k��F��'�����V6َ�tH�Q�\�j	�AS�O�D,e�����X0t�!�F��u�����Ju%U�ML��F��o�3���C�r*c�]�atL��1��#<�֛JL.�kl��NH��&�d�\D]DS�Q����o�$���~�g��P�
��l���TG��&���"�����Ar{U*n����f�Sorx�?���?yR���8QvՄ��n�0��N���U�y�
�s��S�lO��P�릌)�buӉl`o��w��͢���ֆ�T�BI,�N��yO�J�<��Tm*�؟��q��&�lma���L��S�.��N�
E&-)�=��(	�+��G����Q���<�n���+G��Nr��� ;{:��Vj��+�6�<�
�0,�����k��{�y/���R�ş?,���_y�T����Q 2ä�7�(��!�Xz�+Rp`m����-��(�:60:��iI�X$sv=�C凕|�ϷuXD�y�t�e�sq�Ǯk����13�����r��+�e�,#��G���l��~�*�����"'j��$�J�F�%�ii���1t��1nq�Ģ�+���7��6w�,0u��S=�[��%r]ă��A�CL~y�;H;��+G�˛/�מj��b�E���Ȕ^F"�U����_�K!f��|����U�J��=$(�:&w3�\�I�SM�Ԭ��>uU�?�F1Jv�����:�n�������P	K}<�E�7H��e��)�H8�.�~{
�~��1T�0ɳӿ!�aUH�?}հ;�]�]cK�6�0�-Q��_�Q�rV���v���+�_Z%$g����	6����N}���?��>��.��e�;��a��V8��� 9%��@@b^m��%5@i�2�ڹ�:h�FtT*���k}�==�W���"s����I�#�������x�D�������,���	V��/��*�'8����6'R#����P]Cl/F���p6����S�,{����_�W���f��Ye��*d"�.�&ZRD� �㏢.S�J��ke�A%�JkV��*�h�e '��[ c�&Ld)�����ilx9 OϬ2=��ǘ8zz�^�H�'���p��ݠ
�)�y��^�����X��U{J�����������Jw�-�r��EX�1z�|���*��:[~�������D�����)��=_l�$�&��<#/�#�Fч��=t�J�iqqC��QSPN�qIn��=c�'ƊL�g��PR��Zܪ���W��o��A
���XԎ�Y�Ȣʜ�{F/�Q�KB#lx��:�b��Pl8�b.I�̑���E"��@� f3��Ib�u�� y����z�-a1?P3�\���܉��G�2a�����疓�W�t�5Z���n���֕+�� RUy0?��ioJ9�R�&4���&�6%7wA0�y�σ�1�d��		���;ߡǁp����ׄ��v
�"핝{��BU~o[�! �4)� �@�V���ӳ��N���:�i��mtK��>p�ͪ�70�����đ�D�&�����M�|ˌ�/�Qh�͏)�1��bYVύ��q�t�%]�~�Z�)�+�أܣ>*�5��e�|:n(9.�ZH�_�Q&J;�)�2)!�g�0̨2d�K�?]�y��&�Iu
T��j�o��ú�/���2�K���j�����rBa7A����0���Gy1"�ۺ:��gL�ʞQř��sz	hâ�i*Z�aUF��r��r�>K�ÿKF���a���b��M�k�f#M|˘��p�*i�J��v�0�7َv�3p��p֢�ǽZ����h�<��ͷ8��H)��bx���[��Ծ,7�y+:F��u��@����y�o̛"�Bx� ��o!w�������a{j4�?����a�����wp
�x�m��T��]����^�+��ft�?����A���8 � ��V4\��p�!3ѭ>�92:m~� "ǉ�����+����LN�Y�ˑ)�ϧ��]�����m��ZoH��!\�G�ǎ(s}򢷵���w���a�jYՖes1��FEֲ��ّNYI��
nc��7�ƺ��'b�Y�z�ף)-�L���om�0`�MbU��c{v��n��S� �9�q/n�e�*X�3���tw�dcs���ph{ڷ�$�hC��^:S��b�v8%L�\Va�2�y���[ZX���0ޒ<�ycQHR��';���������O���z������,2���!�Pl����-�	�T�B��p�{��{>4pA� i��ā�ߖ�* ��� �d� w	2�~<F�5 ֊�K�Ɨ!Io��M�7����<��2\��U�� ��i�Jѕ
K�|w�Ѐ�K|�4yA���QP*��:9�i�@�{c�ѹ�X{��Y�V������,�oIyr>.���r(weD[�)b=]�?��U\4�t�<��L���1� " U&�
���+����%/��]~�%�� ۱����w��F�MR�Bg�ϕm񾒝M]�����P���0B2���/�p&p���QE��'��-u�/��i�^N��ρ�y.��~�91�ʇbj�U���_>w�) N%��0�{�C��{��Cf^�ǚ��2Yg��ش}^$���43������?'�Q��Y�� oZ���	��d��9�0�a�$H��T}7Pށ�t�%g�	��9gJك/�\.c6����Q��dg��r��N��C�)��,fy݀X��:c��.���pm��]�΀��D�tx���2O8���X�=�*ߝ������t������z�n��j��k�%+A<1	fL[���w�&�\*n�`��Ǎ:�������^k�ңk��!� �1�.sRf"~!�z�N>@�S�(@�nH�s"���PhP�&���2'䎋=4������i��/Hk�%*װ�Qͤ��O�`���Y1�G�MXm��r,H�o'���e�\�!{->����k�Ь�ְR�_����G�C�u)���K���.?ꍠ��S�2�EI����9�nrM�����ƃTk?@e��c�2��G��HB�zDHu��X�ɱ��u�#/9���X��\�b���zrG� ���T�l�n|J	�\ۙ C��z�|El	����+�ӭ`h�af�y5Q�$F)qbӿ!~X$�\+|���4W��o������+j����=±��I_����k�i�EL��U�ROO����l_���6p�]R��S���щ�n�HV#@�vtjn#& ɹ�lC�n���'e6u�b�����m�8�ռ�� t�K(aP�^u�&�?A��g�
q׮G ��3���@7*�5�*f>��UC�ʑ���MP�'����d �
����y�<���D�=e帹�!Jx�@����au?�G7	
l�4 �<rұ�w��a�-v���ٌV����Q3~�b7�~bn��Y�s��^yUB}s,<�[)�d��;~��GA��_|uk��=��k�����ښ���{�|
�r]i0#�xuƭ5jj玹�E���nX�5G��h /��|D��3)��U�;}��Ƅp�1�ћ����W{�V8E�z���T���fF�j��1���4Rx�~΃i�f�q(���w`�S��.��mٝ֬r�$�0(r��c��+�KkG#�����`q�4���p�vt�hZ�})�V%� �;�x��͸��4�߻�.59��E��g�2�����<�H��S�I��Wgӈ�36���am�����<fA��QU�"��iI(4��%�U�00?���_31���_��W���a���	�  ���
W3_�������X�����L����#���p5�3��TR>�ǆ	�v��i��G���p�g��b�i�U�KO�$�d7���/�%fNE�y���~a��'�mҮ�wN���#s��ޙ��R��1����+��Ǔ�Y�qa�W��.�9cC�K��8��_����D�e^;}ᴮ�I0d�Y#��:o����R�FE4�ot��;�l~��K�E��9�N�'�8�c���${�4F�[�&ڷ��k����$D !���Y����s�=��IJs���,��)����H�S��=܂X"8v��dN⻄�5#�$�rX���f� �Ym#��L���] {�snCv�\�=�l�g�B��?���m�E�X"$�X�X�]XX���髒MY㒰������ �҈��c�����ѝ���^k�>���i��!b�� �Zխfp����"�A-[-��ez� è|����|z�S��.6���N�=�\�=�B1�eՌb�p�ǁ)2r�͹Z��<��'F����*E;�rpy��:�v���d�a��0�������Z�Y?T��5S}�:�<���۔�)>Iڋl�N�O7xcsSH�=��O�ZqH����#&B�ª�6��1I�� >��w��@ۜ��z�l���/��׍}���p��fӠ�a�e�+ϡ������(tŷ\�5���v�\����lv�b�\���>���_�8��z�*�oW��1��>2��&]Y����nX������y֛�1��MnU���A][��A<E�C��xCF9��%C��)�jh�#��ld ��W�|#�t�T�ײB��&;��q�),[ ��p<��Q3��k����ج\���$J��l��9ՙIU��YSjU)FA�J�΢T=��%�J~L5�w�=���a�&���R��@�Q$I@�a��4۹��E6?*���v��ժ��c�
l�<�0�
4��Ջb��
:z�T3�����R{����;IB�k�����n����]F���ED7|�`��d��S!V��Hy!g�>W3�k(ڨ`5�\��B���� d�6?
r�(��Fn�*~�|)��]�<ڔ��&�[��`��%����o�iZK^%���n�y��g&���|��ݦ�	�%�$���Wj��A�f�����zf��Iuh
���#L��"4h�HFL��Y��"�g�x��g1�G(��!�p�ZS]`F�GH�%$ͅ^���u�f�I��.��yr��^�˗��k`�u�BN/�]=��U�XǏ�(������\��}b��<���u�3���|$�ճg9�G@�w�W����x���.��0�J�Z��%p��r��y��Z@:�Kyt�i;?��zu�'�j����Ig�� *#tw��:�� �����C�Ea'Z��a�_�L�Oi�'ah�[;�kQJ���/�D�C�^�%Lj�]R���5X����jw���[��'u}<�8b��}R;�PC7K9��(Y*dr�ac�����'���kTA3�wŸ(ju
��� ���?k�	/�K���A��=߀KN��wB����:j�UZ��K��}PE�/���W�W�؉���Zݭ�(�n'�縨\�2�2��z�p����k�7����U�0'��~�3�|f�F��>
%a���A��K�MX}�	O�aS
u�zA���ܿ�#��cT�y���m4Ȕ�+5ʂ�c�QZ:^y�XE��WG�^6�d��9��q�V������w�[�H.�[ ��{��`
�?���/v?@��2	�m�����̰�6vq��w#i�$g�}{�dJi�,2��UU�l��)�3�x�k#����T���G<��;��& ���H�Y
�Ԕ����$����K�3����[�8J$����/���/l0��梇Y�����S���w[[�����N)�^�l�NTrC�}}����'[�U�H���1jL����;�`�|F���i`����iS�lk%I�z�>��;/�)�r�c�FH���R���&"��]�z�B��'<���B�i24�KS�6�6���n����u{Fc�f���2R�9��M�@v�/F���j._��Y]��3�et�.�vԻ����Z��<�G~9<�T�KUrE��� �]KGEC����� 3�A<-gb�&d�d9Ln�����o����yy7y�G�@2;�� &�7|�)WY��(��P
q}���;���ԫ�[�;�o��*��}�:)&�:[Mg9B�8IyH���V^D}�O�,PgsBM�I��2a�)RC�(��l�_)�~�h�Ւ鉍.ed�U�H�M�ǃ.٣��/���{�8
!�(������<`�F@��r���B�0o�e�q�;�ϾG�Q:E��HI+���{V����&A��Ԟ��ż��oC\K�$�/�@��4�jUڳ�;w��7)M6���ļd ��!�a��5�
˟�o�H�4k�t6�󏵂�*e����:�شg�y@2~u`��,���$L¥�����Q0��v�o���U)��J���SD~	H��U��BYEĮ�L��-�ulp�K�1u��pG���ƺ������F��/�t���AA��D���X�n�]X�C�1�)y?��W�Lr�oq����>3�UD�ve�P�Y��$���R���F������g�7�菰�c ֍GcG��Ex[�4>ȐL�^JD��@��S/աx�Z2.�)���It�3��\���u��M0�����A1[�Y��tEql��L��V���/�L
�=&0�\�}k���`m����{$�|��  ���AL&�4�˛��:-�,�hU����a�)����6����<��교�tq0�5�3�
�Z�	+MX�>=Q#�YGÍ:�;����@���N���O�+��6��P�9���0��Nt ���ϩ��4)>i��n�q~�qW�M�'G�f;�O~��]�1��4Z2_l ܄K���Pg��m�xFo7� eZ���T`D�.�����ɮ�3NR0D{5m]��K�=�Ov��j~9���m�Wx���|Sa cUo��,ӊ�s�T�q�*ƐRv�%fL;�Sda�E6�����h��V;��ut�,��p߮㫘�pt&�&0�Qh���,"Y+d��)���B�U�!��r�p:�@ć%ч�w�zX��uH�A~Ob���湔����:%�%��W��0�x��Y d�<�}Hi�Z����ã���)�U��M^��h��Y��F��6Oq��,'�z���/&�/��F�R�٪�V�Q�i;��t�x�@.�*���(RQj�L7�E�v |�������~��k��r��z�#��@S�xV�B������>���2��Ki����Ӄ��">����t�g�U2S��fӨĿE�/0x��B8���0���G����=S��[p�n�Qg��X$S�c,��]du�Vf)����<"���t�H�u�!�o��lH��`9���ep0
��M���<��)���݌�-B����*�֖&�l�;�숤���/���m�?��m��1��H\.y�����9�F,y�2��#���T��UL}3�n�r_0
��}ے��M�nu�M�a�$+<���|���!���v�^î��� ��#�l�gk�𳃦����/\c�嘹���Sw�� �3���5�'����^�?�5�p�«K�A�1Ǚ�!�P��$�I:�L��6������ym�� �����_�`_e���s1Xf_��t	�S^����*ɣ��?���.L�%5;p[ g�+mk��\��gr�3υi��rH��
h�:�!y��E��l�$�I�X@�R�C�YG,�����>�A�|�����y�Ž�XBl������'"|�A* >���H꫷��YU�L��/"(���? �,K9]o�;Y���9�G9V*�W:׫�Oa9�9ԗ�ZW�BL�n$�m�6
5��d���/�2�!d���*�5�M��<��<�8<h��BQ��`B���b����	TE����NA)�$�2ޢn��1;��u��読��G�I�qs}�+�B�5ߡB�H�`+!q�(O)Bd_�s��-����3�/jg��	� ~iyCP��Ӟ:����SV�6N�͠l�?��!�=*.X���;0zjS�n!����*��� ��K�+4�r5���E�3�Y/��p�K��#p�_���M���y� �|4xޑڪ]��qxP�$X6���E!����N��S�\F��]�Ҵ4�wQ��p�U�>�������?>t �T?Bm�x�׮S%;�w����8��ȟp�K{��e��.���4�7�P��b�c�VQvY~�.�MA��t]y��/*r��2U��S������_�%�t�j�wE�JٮB��~�����9d���<�l�l�#���&���FDQ!Zf���iT�щG��jq�1�������0k�{�f��@m#���w�:C�ޖ�֊NՎB���"0��n"��s�s�K1H�o��:,(7������nAERD�63ܽ{O��j� �m"Kk'�㌝�ů�S��V������Ca%G9I�I�b%��R�-!C�l�=�����Q�/��0�w��,E�"��#�J�o)�|�|8� ��B����F��!uA\����f\n��>�83Of��u+Ӻ)8R�[O�O��ˬ>}>iY����Ɉ��A��+������&�m�bRQO!s������.�i��z�y+�wng�2Qr0�RH�R��J������*ܝ1i�f�	���ҋ��k�d�S��S�9M;�q�v�?�ٵe��tb)��v�ϗ����h�?�#<4"]<��As��W�AQ�ٟ��Gg!)%R@�=Fi�J
N_(3��Xf3�3c����d8[5��	����&����n�;&�s��	��.U<#!d~k�a�U�wN�LO�c�\��7�m�#���&hk -x�:U�U���Ijt����8������<����z�o.٤kN�2�c�M�p?�(cR����RyތԳ,��(2��[�;��v�>�pJo���l�iBG��B�Sh9Ú�	״ǆ`.H���� �#���(I�6���]*9��>F,�*��dx�0�s���NLh������w$�$'�rb��j�w�m.w]��F�M�?�|J��͹$P��y3�/g!��S��ö��S�2�P�6�sP�q�?h��[¼7��g�ղ#qZF���]���K�V��w����n�K��Y/B�z�.vy�>�mA�c����a�[��y��cL�4����72o`���C���֢������V��	��&���1�4o�o�b��#�sV�b`62=:������ d���luW:|BKv'l�������v�����I���n�ϼ�&\^��"���A��㪜!�%��f�e�Hɂ
i���zߠ9�:���Q	,�A;k�����3����k�y��#��D6`�����6�:$��BЂG8��l�P��Ņv/����&���ʍ)1;+$�a
�T�h�Jo��>�J����N�Ed��a�tأ�h8�<�ᤶ6l�+���õ��9R�F{%e�!��"�ʽ)c��J�k:�9N�p�[=3Ԗ����ԠY�;���x���7@c�k��On�=W汰�N����ž����"`o�2YR��_�Aq$\H�ڡ����A.�y(�@`�{�o����g�On�Yn�J�fox̹g���'7��+Z�X)��&����e�R����+��v�?�1 ��B�܌���Okf��.�g^Q���O�9tW���]сt�lh����xw ĝ�+*3e����z� V*@���c�ȅ���wWx�&(��4�F��1^'Z��� �ID��=���ߧ�����{/��Z�������k��R���6w�G��8�O�w:x�A�%|��l����#�A�{���r@�1A��`�8_X�k���0Q��H���d�/U;^�<2>���1F��ª�����ԍ�=��Wuw����5��i�\�=��8Za4+	�cJ/��A�}����am���m��i�������]�^�D��/�[�'ox�5���6:� ��"lT2�gGk%������:^i�++l��oK$�7���ܢI����`��}�p�j�3���ш�"���|uzkvc�$O}����ɋq�_0�[����ʜ� (��J(F��]|w-eB2����:fn�b�O/��d����r9HVV_,C���Ĭ��J,��ѣ��s|���5�&��Wfm]d.)�
�{^���Y���\I=�ξ�B��a{�M�5��C�#Oeʥ�=~釻)z��mmC�(]��z޸��I\9����ضy�`;�3�ƞ��]튁?z$G�=(��ޛw����<M��b�r�NP25pۣ����𒞂�Nf'	Ns(pdӀ�p��*VEFt�H�e��0~,�h����P`�mY���C��`�U�N�k5�nJ�zMA��lY:�P���Q�'���5�
��&_{���!�_V6Fe�;���F-���"�
L��&��Q�~���|�tzY�=Z:�%������	3��:R�6D=LnYk�ؖy�n���A����*'�`2�4_c����/������a �B,HD��zHX��^Jt���+}N��\�'>�b���橚���dY�y��ٰ�4"��^f#����p�gzU�c���'i>4͇��P�����!�_�~�&Ux�2?0�|��Zi��tϋH��P65��������UZ,��r�H��?J{��MQ������y�#2��^bV�a�k-,�U>lC�G<���2�q3RJ5�����$i���f�g(�юG R��v�"��dh�}�v#~��O�f���.:��T'v�J�ђ;+���9Tc4��
���c/�h��
�g�LT�B� �g>f:�8p!ȳ�J�>Ē�Rؔ]�T)M�ą����L��B��M9��=R��Fѥ�a4�����L�]�,��M�E��?�%R�" ��5��4	��M\���U��	�q�L>�T�n=�u|f�<;�	��X�X�$�:���ϖz�4�ౡ��g�$.�Y�b/����,�s�o��.��-�'�9�*���\b]�]I�#eB:�Uܩ,��ro��9%� �$���7�f�����*=�8E#�&�)��FW��a�^��V��HXK��!��r#�}Zp"zF��vq�C0�I-�� 5��8���\,��HO'�p/����z��xÖc�)>��}���y�y_$L^�su�,'*�!��l��"�a�*�F���Q7J�_���R�9�'r`��\n�a��rh�Pǘ�fw���#������_�%)��˯���a��S�y@Zt�K磎��G�,��5I��٘��a�=�B��᭄O�i��N�9*`.	�C�P@�y���nW�ǫ��Kl�w�#�x�Rs���t�l��bq�q��b�ΦV'f��]�ht�%Rr8��(��Ȥ{d.�d���q�N%Vi�pڪ���:?��y�,A[�m#�D\�r�~{%���O��il�T�3{X��=����\��@K��I�d�P�k�of�6���z�s.hX��M�l^��b��J�@y[A��=H{䟬���Ԅ�Cϐf;�e?-����<�d���Χ?�ݙq�
ZF�k�t��U���c� ����0����Pő���mB��6f�F# ���i\ 	x��}VG���4�Iw��N/�[UWR����Mn����ed�!�E;��'Ž9�=C>z�v�v �T#{�p&��o��Huk�QW�`GU�ѽ�e�u�[����v�r�p��{�\
��K�#&fִ1�k�?ci77_��"*��/�����M-��*������.�6��t���mm�GHc�4_B�͎C�}�1h#^S�޴�>�CCv�\+B�D����xF�~K���I���~5�m�%��x�J�i�t�Ȳ�c@���L~*[p ��T�n���`㐿h���L��Dʖ���wC3�m��:�&5�%%Pt:t}M�S���G+�C��;!��85�	C���L_B�8Q|�߹�M�h�"�q����y�ޛ<[��^T�H@	�a�sH��ش�kR�7�˲�@_�(�����8ļ��C�(�#X.�Q4����C�]�.�g�d�� �=9P͚NIL^`&P�XƷ[�tJ\�`���Vf��fw1���R�H�o�+SaJu������8�d��ݗc���8p+����f��Vyj�J���M�O��*��a'���7<��Q%��@E�w��u� v�tF����6�7쀏46rr���Ѭ}B�i��d����[��q�&+z	��
4�d]7_t�kꐛ�ge�$(�ķ�by�ϚT���3F������v�i��S���s�V��QCN�Y����J��z��N�_��T�{�l��������8ۉ ��9�F�5鳀BP��Mo�	V~}�`���>�6֐+��tK��l�� .��+]3���Qͦ5���&��$L� ��6{�\�5���+��*�P���X�����o&vi��L:5�w�������`Zj��C� ���oZg�ē��o�li���>�%vC�/phڏ�9V�w�AZ\1s���&M��p�nA��X���cv���P�6g zP`"�ڧNǕ���W�B�?v{��Yݰ��jL�LOm{(y���&���L>���5�޹0��<��rĔm�(��_�6��$2Ϊk���ڇ�؏'��J�zfJb��`�zSA�n���eq�毰�	$�/׼�v���q��g��P�H�]����Ѩ f����qH�O�cs�k-�Z�+�<g��Ӿ*w�$�+K��8�p�Ev�[\X|a��V���;RSy�ٶAk�Q$($�{q�"��q$0���rS�SnL�:�ť�H���vpF�4��N/�O��ǈр���V��'Q9� |c<�D��`.�$�����ؖ'���;�>�Y��'�d|�!�sA�|p�5�GP� �\�P�&�=�՗�d.A����d��I���>Y` wBE��a\%�FKcohJ���[���/_��z��bGb\vR;H�	� 8���v�b')Yj<���y&���'$?���S��jE^%����Ŝ+��{�������Ūƾ��� _*׉k�n���$�9r����F�G/F0F�b�ö��	�7�X��8eYE�^���^�N�r~ꧽg����j��m����Cc��~�yP��<�(�'70RtFO}��ˮB�cZ~�愠 �zEe]����M%�9pm��v��Ș��i�XǤ/�e����XkS�0�����I��|#w�����
�*ِ��4�M��6`�yN��~�p�A���5�r􃢑1f��-��.N�K	�o����mW2Ntg{U��я߁0�g���x�Ȋv�uD�ȑ)�� TD�1/�˺�j���3,p��;���S�	 \)�6�^��%�a�!�c@2���@���nS+f��B2�ƣ�S�Ui�ܚZ�����SғK�z0�o��IZ�۾�F�qt".��mG�����jv���a��<t��"����h�VD�3��3FF0A�oѐ|4�GC^*Q���d� ��j�Xڌ���j�!m����/��\��qo'r�v�]���DA��0��#,��=ѻ�������O�o�޳5�.�i��dN<��3Xz,}����)Z��6L�e��kJ?SO��xǋ���E]5y��ܮ��U/_V��`�"ER #�&I)]� ��=d���[�J]W������?)�h���9����_�I�GuPS����L�;�9�7?'$�"�\@�T���I�l<YO�1G�翃Y��9:�6gK�Ɋ5�� _�����X��:q�B�]A���jV�����76���8�͉a�)Y�đ��[6��z�@�d6�j�]�����w$#JC�:ԪhHr���_w����~5 !."�U/=fUѢ�C:4	���oKf���� A��[�Qc|Yt�F�Y�*�j���_pD��$)b��a�u�� �����w,B>�1G.!�K����~�Lj�dԍe�P�O����Js�ʨ#�ܹ[�8�E�d%�4��M>}MW���bpS�H�j�)�r߁�If�z�qs���ޒ�p�q�\_�]|?��OҟM巷���:���k�%Q,�߅�S�8��
�@�=V����q"WBn�o�Њ.�&��>VذS� 5�غ��SN��m��]�t��n�qJ1L���g
]5@��O���P>��c�_�}�uIݬU�~����ޥ�Ί�B�SZc�4������s����U�4�?�V�,H��p�ګ!�2.��=��Tz夻�N���������E�6�t���k�����h��|�,#��1����ʹa�'�ԫ������.�p����D��.�"�=���b�Aף��k��_�<by{���@5%�t/��u��R���~
yysL�OvX��MӏTK�졩2���,v�0NaR����&j 1r�����~���7��g���e-�44�:��J<��p��|2�
q��H�^������}tE;y���~L/m� 8�`�ƒOk����}Z�D��Nfo��Li�B���`�Z[o�"Hm�M�{���*���=Q���V���p��Ds?�XsxUH;�ek��"�c��Z������ѫ�U؋���G��Ư/�˳ᧇ�'�8���]GS��ցb~$fKá�����и�ȑsjxW�A�vX.��w�������1�9�_�eg��Ǐo�Fx0���@��!;��^U��O�;_㠊�WY�o����y�/	���7jt����)�H<�ų#�ްP���i������g�'�=��'��x�.�H@���>�P[�c"��E�5΄�.{�yeg	�<LN�W��X��͐��I���Zd��#���AF6�K���KP�q���:�U�C^�H�E4���v�C�$�����w�67G@�g���{�r��7Y7�Z�A�v����2pܸ��V��\�]v^��'-¸0h����Ԯ�Teh�v<C�V��CSB�Y`"	+n���x�w��|m����o
�X��;�� i���'�	��Z��`�P{���E��#Dhݦ)W�h�����Σ��uo�^8/����
�,�n��p?4���U�*����"j���x�2Ҩ	��>X��M����-�j�遦[<��PfvX���4���d_�%NM��9o3�~к�81�ҟpEI\&ڨt֎�`��55ߏDs�B���|�Jk/�v��ȸ���<�
�M>��*�s�"1Z���A����ݿ�#�}��h��Q�?)�W����m�L��e�N�t�ajǷ-@�ދ��y#Re��� h֫Cl%@�˨��5�Ӿ66�h��hw�r��]��^���7B��"'�;h�(�d�BO�����̌;(m?8+ =�)��@�daZm�%-9��h�2h5�T۲čQ,<��y���4�Ez��G)������W�.��ނ5Zx����"@y7��M���qS�Vm$����[5�c�R-��L�?~A$vO��*��	6����XŴ}?Cyݭ��n��X�ù�3���r���~����o�ƾh�Rr����3�q�N_7^�P��u4����؅£�&��Θ-�w'�g�0��|n��t`ؠ%�g��+�&\S�}���S`VW�� �7$0!evIe��
)t��uk�c�&g�G�x`�;`\t�u��.aȕ��\�f�>l��,Q��h�'9R�8�'	7���w@�p��g���n8�4G9���=Z�Y�I�y�����Z3��}z�~��,Ӈ�>?%|)����1xKzl�Ea�+)�dt�� 2����+���/��V�<�,�����C$_�\���%gZ�B�B����+"'����gN��;#3��,���ŽI�B39���T�D����G*�2���/1>�W6>@nҎv��6����<��tI�eVt�����8w����A��`�Z|a�oM�X)���u��/P�8 �GJ��v6��W���U�$斷c�����.�$o�Qk��̇��	�7(�>V�_��r߳+�*��<6$+������;-��_t熜v�cH�`���L�"��ǆ��c��e;��7t���C���Ռ���	��z�l�%~b��F�>�����Į�0w�,k`�		XJ���I��DM|��&/ڬ��� �F�H��m��Nu;��t�%�t/�ymU\+y[���o\E�h�y�KbD+��h"��^W��T9�p�����H��F|`--?æ�^�۾&�قqW��Z�Z���>F����-��,�v�\�����J ��qt* �\Z��m���kv{����P�y�<�u!����^y� ���x�ݧ�Ɂ$�]�\d��7݌���,�΋�yt������%|�I�S*�a�����l��L(|+������`����V�7�Ŏ�SkQ U��*�dfo�6�Bo�`w�Ȯ���Wոۤ��*�����`�X�W?�U5M�r�z6�8("�Au�i�[9���I�d���Ź�N��@��O��)�����r �J �G0.�B��c_v��TX�x"u����Z����cĮ��� &Hv!�����^O[���R��H�H."�٫�ʗ�1�}d�/Hpp�NC��=�!^ҏ:�_���0��u��[}�nՄ�hafAC�nԷ�][�M�Oj'E���T��=	K� �A�Ǜ��4 �֊-c�W��?k�/f��W̳�W  %��ܗ�����Չ��P&S0�Q��b���� @��q�yTETj��q�zh�#�~ǖ�y<���J=�k�b�4��)�׬Ev�f��%�)%�ef�t���h���P�<vY�(��O���_�s{�U[���
C����9�o�t�(~��ޜ�s	��,�>"�J�&�K����4}Vd�w�0�FwmOj	X������-\6 i>�U˃P$���"���/�����?CK�֐ի�}�w[/���1�#Ѯ��
���n�ʍ)�n�����B�h̖H-N�gJ���׍U��f����Ywl ��.���6�X��D�U!�7 �E�/�ԝ��a6���Q�Z�=�2����.7�+pT ����%�I��6��i��h8�����
z�a�o��+��Ԓ�f�v(����G<��C����.\�{��ԋO��w����/�kP@��'H��x���!^[��Wy{I������'�`cO+v�[ ����8���w��>Q����'K��w[�@	�4�7OC^@2���	���w������ޗ!$dSF4"��f�0��zilۈ��Wf�
s,u�,��5���fU����>���~�Y�8�xY��[�!��ǁ3�ny�V���q����1����E�\qc��1���	B�'	$L>��QH�Ѿ�o�\f\�����o��z��[��?�ǭ���,��bR�k(�^f�'Qc��Dw��BfW��e͈]�`�[����
Ex��~!��V�(L|tU7�)_E���n�(�.и�3��	X�N� Z��1���K�y���{�\Vb�z �K3��A�C�;z^��{�@��ء�3�����+��Ӝ��A�Yy���h����7f-�PO�A�j"Ih��i�'�fi	�PD�GVHZ�>�'��z�N���,:Hg�d���6#��c��h��xt�0�ߚj������!7�f��ؙ V`W���4��d�{d��ID���"�F�b��*_`��U��Pr`�*���l.z��-{�<Z���2�b��ѹ1b�TZ�0�[M{x�"/l��}�ۜ�z$aG��#k�q�{�U(v?�掁��s@���6ȓ�)�P��
Q%��iNYM瓲���nf��1���� ��z`����h�=��|��x-���ϱ�ʸ��x,��|�Xo��	B/�>��^7t`A�'�I7�>�<�򸳙�����"�pU�<�S�8$m�����f��+eK՝v0�=�l�z����Ɇ~IGTL �@��ds��X*b�?�|����Ĳwu:�I�jk��!V��R��kw��l�t��f��D��ްI\��!U��E����g�5�9)��v����5��#��,[�묙o?
�^�{js���D�LLS�nkw�R��)����6*S�Z�R�P�x6���q��鉮}�]Ro.�c����9�!���wߚ!'����C����]����' k���Ӟf:ܰ4zf��e?5�j�����)�tfd�W��G�=c��+(}K�E�-�W�S��!p���Q�Nh�QJ�9*�����W�g�D<Z[��n���.똾B�2[��Dll�C�b�QE��9
R��O����w^>X�|��%!@|7F�(cCY�n3���D����5J��<u���g;R~C"��k�@N1� ���z��
��b	�-�@fuS�����`��<�iuu�έ�%~��;2_�gswZV����"����N(��R�aԱ,�a|��;���x#B�=��*��Ck�ё9�!'3+Ȃ"B]����Z#ue�a}��-e׶)K����T]��%e���� 4}���Lr���e�d8���,G����_�پ�����+�ƴөt�	ߊKm��ų�'X���}�u�~`��2���3�r�V��HDl�X5������7�P�g�#��}�S����p����
Џx�ۏ������m�	^�15���2' �W.�7���~�Xz��}'Q/RH�u�6�j�sˀ+љ�Ĭa�ʯz���]VY�Axf�qxCY+��{X�b�Ȉ�E_�D\yZ����>`y���fc-=�gDIc��E�0��'�Nٴ�fC9G~54ҏf�f:፹-�1� ��;�{�?C?�q�N�5D��KǞ��X]"*����
'�Uȑ^U\�Vf���J��t%�P��i`�U�N����6{B��N�VDG�0WV�O���ZaOǓT����~��gJ��@�]T�`=[\�P��` s��,���/
�܍m>�_J� N��m�!ĭ�����2J�����M?���)����j!�/յ������{��4�)�����	]�hA;�]D��9A8*��\�F���;�<E�H�jDG,�3�-lEhԔC�n�vݓ�����>:ݍw�n�t�v&U��Fz6P��r��"�`W�q��������k�%+sȹ�bN.@N�a#��`�o�U�P���V�g�R���F������������W�Q�F�!�ȳ?d�271�B��wĶ
68�.�"M���{�*����-���F6�����͊�m�$���9�����!��GJ�$V���J���:�9��-Y��q5I�Ų�{�,?���_�F�=�{+N�aQ�������^�U�K`ո�z0�`\���p�F��'��W�[EU�vH�LI�]>���#K{c�gK`L�u�u��'�|ɟ��L�h���z|�iA"�gd�:fnp��+�9�'�e�6�O&�g�ן�	v&�ʘ	��:����qv�p��4�┳Sꁇ�QJ��D"��
UT�C�5���H��כ/dc��p��~4�A�"����h�����w��I��شG��Mr �q�ܸn�` �@6V�;s�5́K�E�u�`�[s�Y�%���_���7�ʌ��u�⾎�K��܄��������������]׭˧���ė�޵<e�rx5�O�AĢ�A�v��޺>v��Na�{����(Nj�����qtL�~{O����cxv�%��̩��>�
���{�G1��8������&N�4��rm�%�!�@A��}�ͅ:��;(�j�:l������EC���&�d���#\/��T��V�g��p|����x?L��̝��e���7�/�x�����j��wp��T�PfzQ�4bV��R\iAyK�I�qP�5`Oho�zϗҵ2�f�Q#1Ŀ֨��O�벙Ĵ�]���J/��J�A0�b#S���K��ƞ�mM�^>��+�WE��;i�`D��D��4aJ@GK���*��n:�I7�2�4��!$�bB�����a^p om&$'��^(�]߼ߤՕ������A�$o�@�Mn�^��$��($���y��T4�WČ�,���C�2��/��c� p'���)���:��\���b�1�X������s,���0�x�Z�u�(��Gp�D)h�W�X2:G��9p�H{����z/�_k�h��W�;}1��Q�lQ�gxA�sM�:K�b�}��c�*�e���rc��o���5�u-��J��� �»�CCi"H�|��>��޹T�nK2���ݟ~��Ĳ���#�i��;�N�-L��ɤr�t��O.\F���a��;������FE���Ɉ4��g3�u�u(���C�ʛ�z|�7��E���XTAtUh*ۖg��s~%�<(��7}�q�U�,Nx�[Zg���Hs(H��.ƵOp���B�oS�e@�� ���-x�o�RJ��|����R�;�K�i�"����E��
�{�
L�LS�Zҫ3t�˂J�-eZ�`����/ewE�׻Ks�-���7����� ���#��0.>��m���"M1�����ҬI^݋��;+F�	t��<0�mS�?��h�!
�t�]��}�����=�<k��L/�槅G�ȏ��,j�d��-
!�8?��P����������rއ���BL~{dV�a�2~��v�v"!!��G�Fι���t$a���B�:��V�2��9�W׽ht>\�����$ 4PW�{�^�P��g�S_� Jm����^��������Xmʉ��&�eO/6�zypE�N�m�}�ʦn~i�	M�:B�ns|r��{y�!�N{Sc�-�X~|���
5Ho��{�+�7'��b��{)�6�݇���4=���ZG��׏z�_�
�}T'�:���x�X�/�3�3��Ҋ�E����Mn��p@-uM�1eǱ���xlv�"�dr�[�tBT%}��P���S�����4��G�MN�s{���?�M<(�߳��H��������ϒ���wY����|�iy�kuz�c��1�)x��5������>���m�	F(F��}�ã7UtZ/������Xblۣ����X��κt7(���H��F�>���c�K��	[�{��[]��ybn^�@m�S~��o��nn�Js�L�gE�2����f�1�hhh�C�q�w�Nku}�+�Z��?n��7Ǵa�ӤISuU�fQ�4�ن�f�����R͕vr���T@W�}���L�~+��DІߏx���<ޥ��%��G��2S^��TF���r�}4�ה�m�_��	߄*���Q^�DI���R��\k��t�g�XP�z���ԋ�� �	\O�3ހ�4���5(&�N�$�ܩ"8�߂@t��Ӿ/m�ȫ�f�p��U����A=������	�.U E�h����Nh�ȃ��b��2�(e�����Uj���!�0�6�[~���<x�:aG�,�lov�ڴ�6�f����3q+�m� ^?y%iQ���5P�h��K�|���`v�名�%�L��⡢�X���YF��朎x�	m��sL�=���nHr�fM�Z�UD�P�²�(����
�y)D�czE5�=0���P+U����#���yn�7��u�]|İ�� :ᅂ
�_�W��� wo="�lY�}� ��������p2	��q?�$U��3�·F�zÒ�{��5zC�ET��n�\7��5��e8;���|�\ d��SN%����L�K�{��_Oߌ�V�m9xlRo�#��+�6 R��&��2a��Sj^��5=��q���������i�W�!���#�N�wX/��4I��ס;���q�"��G���ӥ�X[\�>6Y����w�ā�&?4_��T	@ҹ�%�]���	=�2�/����Ug�{���X8k�	��l����_q�k޴��Re�@E��Q`宴��@���.#W��U���)v:}�>�������&�A����,���YG���+Ï�����-���ji�&�B(�u׍�4�&S���ܐ��OҬ���U'��&;6#�9��,#�p� ���._4�ݡ�_�)x����OW+R�C��D��% l��E��Ñ�َ�"��S��b�\�wf����<C����]�8�Դ'��k%���������V��ͱ��}���2}b�E�Y���eF�¨�$,8�P�@,�D�%lY�@��VF��|�v8c�i%p����-Poʘ�R��6��������cz��:K9��9�.�<��T�Qc��7�D�#��B��F��`!(�*C;Oz�ɷ=�~��2�/��!�$A�\�J�h�l��-YN}_�1�<WoV�����|��rMC�٧Ll�3y�P�w�{R��r1#���ܴĀ/!}�nc��*{od\u�v.�zOچ��^�@���Ӊ)��,��%N����~�VAJ�m�ɮ#��v�NJ�'NM�L��R�D�����:9+�0i0�ӨS��3���S4��̹�!�%T~|u��o]�p��:)����Ȭ-(+�M��%�f@c��`�	ķ�[�A庆����Rg(.�m���3��Z�H�a�m�7�Q�0�\y��e~�qxE6��&�0b�j�T_g��X	��$	��DL�ppȢ�,�N��D�u)�2��&n��^J��~EY����6��]�VM�ZjH�t����/ �9e��oԬ���_�s�H	8��5^ґS��K[�C���hGG;���� +�~���<�T�Wx�}����9���-�S�b{y��sS��Z����%D���W��@M����!`��T�==yX-��&�א%�n�(�Uq+
HS�b����Q�(��ov������{}�ÞbqLO��ՙY�Ə�74��aJ�n���y
�Ix@n�|�X�BJ�w���'�PLNy�q�&���I�������5y��BY"�l�eA�t�Q6 �w�#v |?�Q��:�u,6 ��VE�!�X��s)��|S� �#�i�١��P�i�g|(Du���epY�ɍ��Rm���7���A/��ɤ����f�e��V��ET6D��hU(��L���JFh�1f{�oy�i�U����K�7���j����t�'���1><�.��*��~3�K�#S]B�dF���C|��h�5�b�X�tr��X6�}VW"(��1ű��X �C�Iη_ ?P�r�	$me�?=Ϳ�Me�ft���p��yF��=�qi��	
+��e�u��f6&a-k9���*�*�h�9�z)�3��o?������5񘇉F���;���Ss�'���7걹�YBD�G<]V_�,��Ms��C��?��@�<Q��gF)�լ�K�W�17,10��~Y�W�S��d��a�<SR�d�a����?����Ö�Z���pk�ۋ{����q�sT]�hx)�']�]Z=ׄ�z-u[��T\�� ~F��`�$��#�B�S?G�%��BL7S�H<j�$t��O�/KTQ�b;��z�.�~i�R�y(�0t1�i�g�o��s��T%��8���މ�U�֮	w�h�{�s>��w