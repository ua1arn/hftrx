��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}־���1N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�<4��ˌ�ň��h����mo����/~.)��3\�R�F*}�c}��uO�������~y��ϼ/U���T���딣0&_���X0���2|	p��rw@	@us�犕/�h����
ۍ���yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪ�`DY��Y�Ǯqh��@eYgA���z�Ś��
��H,7O���u\\�R�F*}!����P�>A.hJ*Aj$}���7�A����А��䬣��x�Mi��Zߧl4���0�?�1~�x�c&	��/v�&����?@��(k��yg��$]B�ʇ8[�r��xmܵs�����G�9*3�-�&�Uxۤ�(���.X?��M���^����S���	;�e���̇���S�����g�R�b��j�V��v�rX.�?�d���&�����;�#�}A���nXZh��\�P��}�"7}����Z���n9$�ܟ
sҖϧ�d�̄\�2��s�RdE�̈́|��S��B B��q�-Z����˞f�C��I�"7���C=�{3t�6�2͵�p����d�ً*��\�w�_�`T%�.��1�3u-�&'��Y_��!G�c�},]7�2���r�N'!�W���I�Р���Ӫ�ҋ��R��@2f�)��"ƴ�zI@�ôւ�Ѓ0��K_�0�� ֽRNc�۩<�r�^��	���w6;i����Uͬ@EH�̏�؊�"�D��_���������b�Aկ����<��,�4��>�����F�.�x�w?�f��i�:`�+Pa¡����~������ H#p�x^�4զ3�0�j���d�k��"���\S����(���G=���q�?_������
=��8�z� :����H�%����;i�z�A��Q�V�O?�Sկ�S8a�bYh�j�w��a�[�?Q6H�͑ԫ�N���j��V��jѭ�5�Ϡ��)�NUD60L�{U�����t�1��6H`���ԅ|6ٮ�(�Z�4�� [�_�wy6)qh�x^�`	ַ��K�&�a��|����W�%�э�U��b����=N�C�� c��(�U�q�4�����{U�����)���0Z	�5}�9`	ַ�=�?��3�r������z� 40 ��ٱΥϐ%�i� ���������|�;�Ojz�`�v�e�~a��V�̥�
یfz;Vr�'K�Ē�Zq"�{U�����YI�šCUg/.�3lC�)�Tr�>b�LMǓߥFS oe$�{�$�ħv_��Jr`�F=^�~	�5w/� f4\���d�kⲰ 1'����
�j�GR���%��|$�����6P�������"����g��%a<��As�Gw�b������>�;m���T��bz��F��*`nԡшt��z�����Q�J霝C�C�~�0�
n�f�)^��ʆIf�ЯmMǮv����UrZ�q�PO40k7�=\�]Q��h���Ѳ��;����J�Y�:���."�`k�0�N���K��/9���-贅����	^��������������`��s
�C�{�(+;���%kr�]Ɔ�	y{�m BM���7r�S�~Di1�(��bX���A@�r$��_X�=m2J�,QZM��2*����v�v���AB]�@�Ț�}�����ʟ6s�zh��/�܄^��R�8�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�sQ��X�zȣc��- ��Ckӏ�^!�:�_c�~:i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�6A�7Oq��@���,������0��D��L���_�L�3��0I}.��dPc)y��dÂ��t�iZ]XF�IV��
�Q@���k��"�,�>E��ʆ�In��t��Q�]��-P�vȜ�[��CC��E\!��-IÙ=�H*.�PS�����k�5l�S2p�Մ�A( ����_ֲ��mŹ�[�g�DPp㧥���*�W���g�JHn��z���z�O҈��O���Ch<Q��T3�F�i�6�Ặ��Ϊ��p8/��e>����C�z¡��h�'f R!�`�(i3N�By3��<�]�!����M[��ǢR�����!�`�(i3v�ј�"��Z鎬����A��:6])2�����Vc2�����Vc߶�z7��Zr
�0�M�yObFT+V��퇇М1!�`�(i3N�By3��<�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��q�\E��0/s�1��p�E����F��j���0z�cUL��`��`�ю�������[��CC�z���a���ł�!r�dN�<@Iv��nt=:�:E��]��8|�;�Ojz���)e����|g�Y�'���Xw&�<���8�t��]�'�ʪ%��1c��Et��q���U�[��N�������lO�LYw9���TD��ό���.�:)!�1%�@�	^���y�E����F��j���0z�cUL�I��6���T�\ ��֕ߝԀ�2�����Vc2�����Vc�i�T� 둨t0����/��͈�N�˵q�׏�T#�3�["���N�DNl��Oh !6�e.��xu	�>��l%i�-��+g^l�>&S�XQ����&`���I��w��,>����C�x�j؀O��_���RQ�
Yl���#�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��^	QW�Q!r�fN�ї��q]�07G#+�Ǘ0z�cUL��`��`�ю�������[��CC�z���a�R�wX��^	QW�Q!r�{F��#��':E��7G#+�Ǘ0z�cUL�I��6���T�\ ��oR��m��%�э�:�rQRт�����
L'���Xw�.aX�bAKj�V��v� ����⎕�(�
t�������2%=dϖ�i�!�B����� j���tN2s��/~.)��3\�R�F*}�c}��uO����������Hp�$-iu�`���`�+N��?���&���#�{�0;�}����\�w�Y��k��ı���$��������p侢����GB<[�(i�$��Xo��/�b�P	ܷ�4D�P����Z�zL͊�q��C.W26K�~�J�� m���"u����(�ґ��:����0@ȹ��ZBi�mR�5*%ol�ħ���$G�0�M�o�Z��&R��(Z�,��F��>v*�6i��
�L�Л�ޢ�-�ռH�p0���-q+�"�,�>E��1|�!��3��zl����b!��uፁ$�������_j���M"��q����Oއ�?t},�׉é[�=�5x�C��6�g�����w0�7s�9���o>��l%i�-����n9의�z��l (�?qE��w��Q]� _ό���.�}�
�?�;�j���Љ����yзq8�Ј'���Xw���,Dߔ��� @9m����1"�,�>E���]�!����w�Հ�>Vۉ�!=�?��3�����3��7s�9���o��S8�P?_������`y���h}Nw���v)5�Fo���'(����1�U���]�!����w�Հ�>Vۉ�!�K�&�a�� ��$��7s�9���o>��l%i�-��B�D�F �%�э��8�>�}���Q]� _ό���.�}�
�?�x�j؀O��`�����зq8�Ј'���Xw���,D�v)5�Fo�",oMG~�����㞣��]�!����w�Հ�>Vۉ�!����0��Gh4M&Y<17s�9���o>��l%i�-5�e`��9�iK�D�b=G�6�!~���Q]� _ό���.�}�
�?��(R\֎u�=7�7K�P�	}p��'���Xw���,D�H�p0�����dܟz$��R�lD�]�!����w�Հ����(S�s�{��ҽ�!�`�(i37s�9���o�jƓ�[b!��u��}��u@:!�`�(i3!�`�(i3�d�٣��c�A�L'�����CyW�f�tR�wX��}�
�?����'�u�.�k� ��!�`�(i37s�9���o��S8��y�)xʔ���6��	���`y����@����gG��ݿ�[�7�C,�2�!�`�(i3�n`5�fK�\w��0]b!��u��X%�;���|�W��!�`�(i3�d�٣���N N�S��E �����6�^�!�`�(i3�E����FZ鎬������_�,��T:���V�����a)��s�}���+�J��Y�{'%s�Ǹ2���;�¬pX��g��U-�e,%�0g����s��&�},fcXy��q;�E�`JcUзq8�Ј'���Xw���,D|�|��f3��X���&R.�k� ����Q]� _ό���.�}�
�?�\���>�s{�%W3Y��P47s�9���o>��l%i�-E�!Up-i��e�����!^���+�b"�,�>E���]�!����w�Հ��s��&�},fcXy��q;;��z�:;зq8�Ј'���Xw���,DU�m#j[��NۥUn�e���b���Q]� _�rs�i�76b�*ҒT"h�p����t%��zxa(􆿳���2����.��DP֞ �'��L��r>�[I��:�E����FZ鎬�������(���:���U��^"4/���°������R�wX��}�
�?�{U������0�X:�r[3Y��P47s�9���o��S8�:��Q�Z��"u��������f�՜�T�\ ��i3�|)sՀ]^U�*�!�>E-�N8�{�����U�4��X�uʡBs=�b!��u�E@.SWp���!�}<*k`Ë��A( ����_ُW$��]^U�*�!��xѴ��zigzA=v)U�4��X�uʡBs=�b!��u�w� �O[s���?8�F�!�`�(i3�d�٣��c�A�L' ��a���R�wX��}�
�?��P�z�1�rݓ�r���!�`�(i37s�9���o>��l%i�-�s��d�\��ʅ�-`�߬�F�<�;z�Ni��a��*�0ޑw/s�!g#T���Ӫ!�F�!��c܊�+g^l���b��M�E�`JcU�q9+t�}��V9{)=�?��3�M����*���ic)�̩ƍ2���lĆJ�g�*�~���J�a$�Y L���}�x"S�#�doR��m��%�э�X6و�cµ�cl�j���b+}y[��+g^l��~��w3*)���!��K�VSƅ��	^���y�n���/l����J�`�B� �1�Á�a�[�g�DPp�zO;_�bZ��C�Y4�1�Á�a�[�g�DPp�$�������_j����ۈnp��5��aki�:`�+P+鍎���+����$��r����!�`�(i3!�`�(i3t�R!ME�em�B0�B��͵h.��3߬���R83��V��	��y��"�0)���Ih�	�;�b���di������A�+�2��h��G�@�/����t�h��W+��W�7�`K~��CĀ/�h�L~��al�N� ������0j|�~{b62�tstJ��:����\o�LCd�!1v!���'���I���P"G�wk�=5���&4 :��	��o����׋��`y���������y�(����<m��v�)y�Eh�ѮYțȠ��ղ]��nF��kJ2������n�͖�������b�Bϱ���"u��������qa�.�����?�^"4/���L�sPkX��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3w�HjW��ǟ,����In�h�u׆\���>��S&Q�f���fa����xy�ˉSbT��;�k
��R/�fcXy��q;If�b��_�1����!�`�(i3!�`�(i3!�`�(i3��%>%��?V��j�c������n�J>U.@��W�6?��u�#�$IX~���~��p�
�t�^D���=����t0]��2�O2�*�����ϸ�"^�j�h�5��
�YW�S7�.���GX y!�`�(i3!�`�(i3!�`�(i3!�`�(i3im�x�����Z���ot5^ݿ牴)e���Ô+;��2ќs\5 ����.��?��wO��Н�:���M��:�j��G慧1���~!�`�(i3!�`�(i3]q>�A�	?\�z?Xk�V��	��y�y�^	#�0��`�7�`K~���N� -5���$�a�Y��ČS�Kq%��M�Vr���J��:����\o�LCd�!1v!���'���I���P"G�wk�١��	;q��QE|��o\U|~���O���8���/�ݾ�9J�c(&�L�⃓a���8�#���n@#('�cH� ��'��L��:�<�zU��AԢ�a\蟦�V_���07��i:����Lͷw����y�<KX�+�#�W��	��hH�1���~!�`�(i3!�`�(i3پ[���-[�g�DPp�⃓a���80�iN�
_�Ƞ��ղ]��nF��kJ2������n䂸�u�,4	���k$ !�`�(i3!�`�(i3S`�@�p����nZY�J�݃�,A2wKaC�IX0F�MV�ҁGG�K�BN
\�[�����:Fa�7���[�؟�-Y�J�݃�,�uR�:l��;�jmT�#�U���e��d9=���u��r���2��}���'��L��˰M{�?I�my$�N��o�/���;
�:qEpk+Q�h'�Ȝx�5W ��̫(� h�ҩ��H�����K�&�a��J�,���{pe�h��(R\֎u��w�`L�"V̏P���-����!�`�(i3Q� �_tt�� ���$�dN�<@Iv��nt=:�,^g����'��L��\�b�a!�`�(i3i�Q����%�э��5)��Z^�d��-��!T��6�F���N�DNlvr5�Dѯ�3b������'��L��d��qc��$)�~�LS�&Kvmc1tSjv�!�`�(i3{U����ơ_�;+�}{U������O(� ���}Dq�f��߆�p�h�}G[���#���n�W�G��!1tSjv�!�`�(i3{U����ơ_�;+�}�{_8�Y��=�}�Vݨ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Fr��ja�������J±�.�Y�ٔ���.�g3Z�)V��B�1K�8��>L�� 9��/��J�g�*a���Ri�:`�+P~��'v�fm�oH�	^���yU"�
hYY����T,�R�W�u�<�h��N�M܍�?{����ҟw�����M���9���ә�MFڸ�>P���U��s �����$�������_j��������M�y'{w#/ B!�`�(i3!�`�(i3V[B�5�m(@X~�H:�vE��=���Y�_-]��U��)���}�%���4��N�DNl�Ttσ�;�����g��u��D1!�`�(i3!�`�(i3!�`�(i3!�`�(i3��v�)y�E��+�R�n��^(C<�ɷ.7�!��c�r%�ƨ���^R!�`�(i3!�`�(i3!�`�(i3!�`�(i3:)!�1%�@�	^���y �A���EdS�|���(R\֎u�C�Gυ�B!�`�(i3!�`�(i3!�`�(i3!�`�(i3�r���h�0��X���&R�m&�'����X���&R��p���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�\�2��s���1�, �D��u�Qѻ��X���&RWql���,(e�%�<{y����i�q,?5q�A��x�+ż٧��jd�C���m�ڨ�hծ8�w��U��(R\֎u��8���Q�ݚ�Н��ݗƩӤҳ����`!�`�(i3�k��M�KK�+��o�Ƀ�?PA@?N�&�bM?��y�!�`�(i3���̰�!��U`�PW}D��ɍ��Wsp[��X��=@'ѥ���'T���+�%�э�X6و�cµ�p�ֳ�맅2�w����:��q�!�`�(i3�\�2��s������x~>S^Գ3���ƍ2���l�!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��՝� s�#���k$ ��'T���+�%�э��8�>�}�k���������|e"��'T���+�%�э�X6و�cµ���(A�,"T�z�D�R!�`�(i3����H��X���&RWql���j�֎��5s�FF�?g�j�P�&Cd�c����O�*f{�k�(Fj�V��vi$'�vu������&G!�`�(i3ݑ���&�d��ҟw����f�\%M�m���!�`�(i3��F���K�&�a��i
�i�w״$(�>g�!�`�(i3��w�w:�!�`�(i3��l�^!Fڸ�>P��=����h���}�%Dܭ��}Dq�f�!�`�(i3�\�2��s������x~>�"ª�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3)�{6�U��(*�O�q�$��]Y!�`�(i3�k��M�KK�+��o�Ƀ�?PA@?N�&�bM?��y�!�`�(i3���̰�!��U`�PW}D��ɍ��Wsp[��X��=@'ѥ���'T���+�%�э�X6و�cµ�p�ֳ�맅2�w����:��q�!�`�(i3�\�2��s������x~>S^Գ3���ƍ2���l�!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��՝� s�#���k$ ��'T���+�%�э�X6و�cµ���(A�,"T�z�D�R!�`�(i3�\�2��s�(7�Q�S^Գ3���ƍ2���l�!�`�(i3D"ۡ�
",oMG~�>y�pA����v[v%��%�э��XW�G�<b~*��s���v�)y�Eh�ѮYț��N�����1tSjv�!�`�(i3Y9u��4 :��	��7=-�ˣR31tSjv�!�`�(i3ݑ���&�d��ҟw����f�\%�<4�sg�!�`�(i3՝� s�#���k$ !�`�(i3(@X~�H:��}�S�74/������SY|d!�`�(i3HN��R��bP�63Z�t!�`�(i3��+g^l���b��M�-��h��ƍ2���l�!�`�(i3UI������%�э��XW�G�<b~*��s�x�j؀O��w���B}�����z��5s�FF'l/7w|]�o
�Z��k�G8ګ!�`�(i3�A!���j�V��veK�	�$Vͬ�J�������n�0R��#���n�zq������2+m���Js�;���!�|D#o�]�ʄǘ9��V�9!�`�(i3�$�������_j���"{Q��J ����:N!�`�(i3T#�3�["�Yr/r��� �.J�>�u"����!�`�(i3�_��>νrj�V��vG�?-�D� ��U�_:��}Dq�f�!�`�(i3�\�2��s������x~>S^Գ3���ƍ2���l�!�`�(i31���~!�`�(i3(@X~�H:��}�S�74/���@�k�F��w!�`�(i3T#�3�["���'(��Cw�Hm�̊��NM���!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�G�&ց�*�
`���n��ݚ�Н�T#�3�["���'(��Cw�Hm�������z!�`�(i3�եH��^@9m����1�'����u��r��!�`�(i3�$�������_j�����ur�?lqG�kk�!�`�(i3T#�3�["�Yr/r��� �.J�>L���}�9�C�s�4!�`�(i3^	QW�Q!r�\1^O� �Xz���n��뾦�!�`�(i3�����!�`�(i3cک*�;��%�э��XW�G�<b~*��s�x�j؀O��w���B}�����z��5s�FF'l/7w|]�o
�Z��k�G8ګ!�`�(i3�A!���j�V��veK�	�$Vͬ�J�������n�0R��#���n�zq������2+m���Js�;���!�|D#o�]�ʄǘ9��V�9!�`�(i3�$�������_j���"{Q��J ����:N!�`�(i3T#�3�["�Yr/r��� �.J�>�u"����!�`�(i3�_��>νrj�V��vG�?-�D� ��U�_:��}Dq�f�՝� s�#���k$ !�`�(i3�(R\֎u��w�`L�h��=��޵����yr�!�`�(i3^	QW�Q!r�{F��#��g�+C��sJ�A7���ݚ�Н���'T���+�%�э��8�>�}�k���������|e"
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н�t�td���5G�&ց�*��JY����VA�ڦ�c4KK�+��o�Ƀ�?PA@?N�&�bM?��y�!�`�(i3���̰�!��U`�PW}D��ɍ��Wsp[��X��=@'ѥ���'T���+�%�э�X6و�cµ�p�ֳ�맅2�w����:��q�!�`�(i3�\�2��s������x~>S^Գ3���ƍ2���l�!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��՝� s�#���k$ ��'T���+�%�э�X6و�cµ���(A�,"T�z�D�R!�`�(i3D"ۡ�
",oMG~�>y�pA���(4G��>�0]��2�O2�.+��W�
�@�����\�2��s��W��7=G��Hb� h�ҩ�!�`�(i3�(R\֎u��w�`L�y���;�U�q��ڍ!�`�(i3x�j؀O��%c5#	�.�X��ͷ(�-���|e"!�`�(i3x�j؀O��(�\G�@�L ����7����|e"
�:qEp���,��\����0��G���_��b~*��s�x�j؀O��)����bX�'����u��r��!�`�(i3�%t̓�@���{
Bk	䶙%T7u��2�!�`�(i3^	QW�Q!r�����g��Mt�꾸b+}y[!�`�(i3^	QW�Q!r�\1^O���Mt�꾸b+}y[!�`�(i3�����!�`�(i3ݑ���&�d��ҟw����f�\%�a�݌3)�!�`�(i3�_��>νrj�V��v��=����%��v��!�`�(i3�_��>νrj�V��vG�?-�Dn��뾦�!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN!�`�(i3�ݚ�Н��ݗƩ�J��n���C!�`�(i3��+g^l���b��M�-��h��ƍ2���lĮ_��>νrj�V��vG�?-�D%��v��!�`�(i3l�L�`v��A�qIp��KΆ�������-����!�`�(i3�%t̓�@���{
Be���C���������ݚ�Н���F��=�?��3�����3��K�VSƅ��	^���y��}Dq�f��	��x��ݚ�Н�ݑ���&�d��ҟw���Z9�+	҇	��*��O`�� \)��'T���+�%�э�X6و�cµ���(A�,"T�z�D�R���%>�rGO�D mWN�ݓ�W���	�N�M��/�9ސt��+�t2�4��A妡��M/*�3���X�zK;��t��:!�`�(i3�\�2��s������x~>S^Գ3���ƍ2���lĮ_��>νrj�V��vG�?-�D� ��U�_:��}Dq�f�^	QW�Q!r�{F��#��g�+C��sU_GD��W�ݚ�Н�t�td���5?�{�X�[�g�DPp���ܐ�}��ZaEUԾ�� Uv@C�
]�vp��:I�#��u�#�$IX�؝��^=�'�,A��89��A$�P��O�@י����z��q�`���φ��<�6�3�;5 M�|#HK�����qD��=a�^7�1tSjv�?V��j�c<o�;)�yԌ	�����e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�_��*��jC��6�g�� ��-O$U1tSjv��wӨj]h�u�#�$IX���O���{U�����q��Ɨsfĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxV�/e�,���NۥUn��O��\�EOJ�uxmNۥUn�W��is�φ��<�6�@a� ����C�'�ąC>��Ӛ��S�J\7r��*�t�>��G���\���F�`y������T�8k��.ͥ�H�RtV�^Q� �_tt��`���`��{RT7b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3���ըR��Bft>��G��Hb� h�ҩ�?V��j�c<o�;)�y�7u�T�M#d�c�r%�W���b�0�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�#Jh�m"3��`���`�(JŢ��EOJ�uxmNۥUn�Wql���t�p\Z|�'��L���m�kb㳒-??��$ō�Zm\ާ�����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3�c�r%�Dbg�E�%���;_��8W�w��fD.W�G�5�E��3N�nS�(R\֎u���y�l��φ��<�6�@a� ����C�'�ąd�G}%����3f��gmJ/���'ž1�|��P�:k& ��-�������̰�!v��� ��	��*�����zNc5�tiND�S���/9�=eSe.��a��o���H�RtV�^�K�&�a�74/����$�������_j���?\�z?Xk�:䩒=]'�Fr��j�W���Y�c��r�Ch��gb8���SY�N��&Y��V��ht��R����A$�P��O�@יߌ��omq�:Fa�7�����PϾ���"sS<GYqcHTX�';��#j�������%�э���'|F�{_8�Y��=�}�Vݨ!��"� +}04~B3��������h��`�����y_�mS8<�n�|#HK��|<��r�*A�P+�u<_�mS8<�n�ݚ�Н�x�j؀O��_���RQ�
 ,��rQ�/m>8Φ����S/�rHN��R��bP�63Z�t�5ߧE4��Fr��j���_J��`U�a�(��%���a���ŕpO"-�R;A�B�H {��u��]'\gWg��	�Z�kfcj��r���(&�L��'ž1�|��P�:k& ��-����^	QW�Q!r|�;�Ojz�!��_�*9 ��b+}y[��=�$�� �e�d��LaX��T.��b+}y[��=�$�� �e�d��]�
�D`�R��b+}y[�w(��,Z��6�^�!�`�(i3%��v�ڹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&G��F������0��Gd�~{�������<>&S�XQ�����FX��N��W��fcXy��q;t} ׅΦ2��h��M��:�j��fZ���oР�(�V��M��:�j���y�����e�����[BC˜}1��}Dq�f��>���5���ٜ�]A����2�2��8��Ս��Jk���}�	76�&�� Ӗ�t$�)�vx�h�C�s�)j�V��v�xp�"�/x�j؀O��w���B}Y�4��1nzmv#.0H3φ��<�6�@a� ����C�'�ąd=��¾ȼ\���F�`y������T�8k��.ͥ�H�RtV�^�\�2��s�5irAz.l%��v�ڹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&G��F���K�&�a�W�^�|���\�2��s������x~>���zNc5��;�P�t�5�׹��L<C%`_�8��U��)���Y;e�iK-pm!9�>��n4s1��7�癆cgR������������ h�ҩ�x�j؀O��`������q9+t�}����@|��璓�c�������t �[l;M?��yЮ_��>νrj�V��v�k�n�=�x�j؀O��(�\G�@�LW���b�0��5ߧE4��Fr��ja�U�ے
��+g^l���v�Z����Z��R��'(��)f�.����j�V��v}�0���b��%�э��h�Gd���{x��O>\ٿ�6�P]M\I��A$�P��O�@יߌ��omq��.��|ȃ����qD��=a�^7�1tSjv�T#�3�["�Yr/r���"���t�\T�z�D�R�Ro�G/]%�z�-uͺ�s�η3G��Hb� h�ҩ�x�j؀O��u�>����?�4V�I�{F��#�A�Pz>ShR}�	76�&�� Ӗ�t$�)�vx��9)i�F�
�oz˸�uK�5��)��z<�ov#��z7�Qu�	�'T8�	m�w���i���Z��hs����ƚj5?�ޘ�JeW{o\��6�o8:4�I���c�90Mj�dL�d�G}%����3fk��{`.~��j5?�ޘ�зBQcCs���"sS<GYqcHTX�';��#j�ݚ�Н�x�j؀O��{dOCe�@�l��p�xB�my$�N��o�/���;�Ra])n#�璓�c�������t �[l;M?��y�!�`�(i3���ըR��Hk��k�z\a��o���H�RtV�^^	QW�Q!r�fN�ї�;m*�z߶{U������0�X:�r[3Y��P4��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�kv޶Gl��&Y��V�aT��3G?�d���&��#}�{�UA�o���cBI��YD�(�^*Ǟg61 ����������OXVĒ�/YK˫�z���AZ���d���!iT#�3�["����:�ͅR]<�YK7͍��|��W&":��;_��8W�w��fD0�ݖ�_J2�H��#�DKIͰ�ʮ�X��:���t�T��?E-h���U���e��_	�Ƽ��S�J\7r��*�t�>��G���xjzӝ���w3��׍�&�U��f��2��}��3�|* ���dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ��;�%�R���p[nۈ�'����u��r��q�\E��0Cw�Hm����+�T[nHN��R��bP�63Z�t�5ߧE4��Fr��jO.�x����n�b����!�#"������X�ƫ��J��ۍb�o��_�Rv�䩲$����E)e|A��`���φ��<�6�3�;5 M�7�癆cgR������������ h�ҩ΅��'�u�i7�����-�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H����|��sQ�G����)�
�M?��y�!�`�(i3�}��u@:(C�d)խ$��+Ut������F��O�}�	76�&�� Ӗ�t$�)�vxV�/e�,���:W��;k<A��݊��zO�\l��=���
%J���E[ˮ�N���X%�;���CxՒ����F*�L��!�`�(i3!�`�(i3�2��}�������}�xc�n��`��X���&RWql���#GOӻ�����)e����m�kb㳒-??��$��Z���F*�L��!�`�(i3!�`�(i3!�`�(i3��=�$�� �e�d��#;�xw��!�`�(i3!�`�(i3��ԡ6���w��B�j74/�����h{���k���!�|D���B�����X���&R�Y/wp�j�V��v
���=b?BXO�G�|��c��@��Y?;�?���	�F�S� `��e�����D9}�Ye����������8M�\�2��s���1�, ������!�`�(i3!�`�(i3!�`�(i3�#�-�p��F�z�n�ƫ�}<��\�2��s����a�v�ï02�okc��;�4�z!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(R\֎u�,��7-u��5�l��Xy|�W�4�u_m�!�`�(i3!�`�(i3!�`�(i3��+�t2��iK�D�b=��L4���w�_n$�%2���8p�X�`�ƶDk����(&�L����$�N}�+c�FP_4��8���Q/�"����	�bV�̗�″*�NZ!�`�(i3!�`�(i3�,�U�Y��4�����0���꺰���̰�!�Xy|�WCw�Hm��/��kOT?V��j�cC��6�g������;q�z_n�ԁD�k���?9�d�Py��D��Lh�V6_����;�jmT�#�(R\֎u�,��7-� �9�!�Q��s�s�{��ҽ��d9=���u��r���2��}�����U��f���0z8#һ����~���U���O@���zxC5�h3]�< :�՝� s�#���k$ ?V��j�cC��6�g��3��	cA霯}Dq�f���Ě�����}Dq�f���M2�}'p5���s)P<�ܓ�Yʁ���Mյ��.WQ��>�����!�`�(i3���y��lD���qt/��n|s�)>^t�a؜Μׇӭ���H��������0��G��e�������m�"TeJZ�D��Jsȸ�"rRݑ���&�d�����l9�̪=���z_n�ԁׇӭ�щRa])n#ݨN��gg!�`�(i3�(R\֎u�=7�7K�P#�+#��]������!�`�(i3�5ߧE4��!�`�(i3�K�&�a������kO�q9+t�}!�`�(i3}�֙Z��K�16�
���N�p4��ݚ�Н��{�K0�>&S�XQ�E�P��U��b~*��s�!*Ĭ����a%��w�ݚ�Н�EOJ�uxm�}�Z��y�&TL�b��!�`�(i36S� �*���8�� ��V���ޕe`�!��:��w�w:�!�`�(i3��M2χ����a�)P<�ܓ�Y
�:qEp�;�P�t�5�wӨj]h���z��l .+�N�R��C����0��P�R�ӚE�;tɓ�����~��$�� �q/r%Ke���=R
i�c�r���M2�}'p5���s)P<�ܓ�Yʁ���Mյ�ё'�{>�����!�`�(i3���y��lD���qt/�����������q�E���r����,�˳�*CyP��C��?�T'����M?��y�!�`�(i3��M2ϼI�)�ݳ��"��ӌ�r՝� s�#���k$ ?V��j�cC��6�g���q9+t�}�ݚ�Н����F��O��ݚ�Н���B/�w���B}/�%�� ;̃Va�ir��_~s�8	0X��f*������&G!�`�(i3;�j����E�
 �՛yS�RD���y��lD��{���4bz��26��*��;�ݚ�Н����g!h!j�V��veK�	�$V�#o�]�ʄ�	]�k��,���^���'ƃ�3�Y1tSjv�!�`�(i3�(R\֎u�=7�7K�P�"ª�����}Dq�f��	��x��ݚ�Н�ݑ���&�d�����l9�̪=���"��ӌ�r!�`�(i3�5ߧE4��!�`�(i31���~�wӨj]h���z��l dG�B3���%��v��!�`�(i3�%t̓�@��܋�n焞 ����7����|e"$f��_Ub�F�S�1 �EOJ�uxm�Bft>��%��v�ڵݓ�W���$ �3�Ϲ��[� !�`�(i3!�`�(i3���:A���@!�ʂ�����%�E�����l����)/^�蜬�^���'ƃ�3�Y1tSjv�����l��}��>�u��M��:�j�7t��'��cN�0����y'�10`��#	�	bt>'��B��)7E6�D�xW!�`�(i3�_��*��j�,����I����2�H�RtV�^!޹������K�&�a������kO'�^�����ݚ�Н�-^"+�K�;��z��l �"�Mg�ƍ2���l�!�`�(i3��M2�}'p5���s)P<�ܓ�Y!�`�(i3ъ�G�^J
!�`�(i3��l�^!ЙMǿI?��6�a��)P<�ܓ�Y!�`�(i3?V��j�cC��6�g���8���$��}Dq�f�!�`�(i3ns0mWw���B}/�%�� ;̃Va�ir��_~s�8	0X��f*�x{^4��*m!�`�(i3!�`�(i3|��sQ�G����7E����NM���!�`�(i3��w�w:�!�`�(i3!�`�(i3|��sQ�G����7E�/��kOT!�`�(i3$f��_Ub�F�S�1 �
�:qEp�;�P�t�5!�`�(i3t�td���5՝� s�#ͅ�簔[���i\�6R�$�R�IT��Xrnz���+�t2��iK�D�b=G�6�!~�%��v��!�`�(i3q�\E��0T����q9+t�}�ݚ�Н��H����fD��j��ه,��7-� �9�!�Q��s�s�{��ҽې���xQ�1tSjv�!�`�(i3EOJ�uxm�}�Z��yn��뾦�!�`�(i3�	��x��ݚ�Н��wӨj]h���z��l �"�Mg�ƍ2���l�!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f�q�\E��0ÿ�����n��뾦�!�`�(i31���~��+�t2��iK�D�b=G�6�!~�n��뾦�!�`�(i3���#�cQfcXy��q;�˹�+�[�G���K�ݚ�Н�?V��j�cC��6�g���8���$��}Dq�f��	��x��ݚ�Н�i|�rBY�",oMG~�Յ$�O&�#o�]�ʄ�< �SS@�
�رjwc�';��#j�ݚ�Н�?V��j�cC��6�g���⍇�����}Dq�f��	��x��ݚ�Н�?V��j�cC��6�g���8���$��}Dq�f�HN��R��bP�63Z�t���%>�rGO�D mWN!�`�(i3|��sQ�G�HOW�[�/��kOT�wӨj]h���z��l �"�Mg�ƍ2���l�HN��R��bP�63Z�t���'��@�my$�N��ݚ�Н��(R\֎u�=7�7K�P�"ª�����}Dq�f���M2�M�;Ss]�k���������|e"EOJ�uxm�}�Z��y��ic)�̩ƍ2���l�q�\E��0T����I����~u/��kOTAL(�z��?�t�ϗφ��<�6��A���A��Q\�_q���i���x��!ӹx�!�T�+��)ެS��B�02�ok�nS����bK��:z6&����(Aw�,��~��A���A3�p��(�g���S�
��R/�fcXy��q;If�b����|YOF@�*���k� ��$J�L�l:�
d�P}4q����!�`�(i3!�`�(i3��b+}y[�X%�;���X�c��J=S��4AL���q�n�7�����%�#�"_����k��J�fc$��b��X���&R�S���4����E���	]�k��,���^���'ƃ�3�Y�ݚ�Н�!�`�(i3V[B�5�m�Z���������P}�H {��u��]'\gWg��	�Z�kfcj��r���(&�L��'ž1�|��P�:k& ��-�������c0zQu�c���i�L����;q��b+}y[�k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�cک*�;��%�э��5)��Z^�d��-��!T��6�F���N�DNl��zI
��Z���Ӗ���7���U�� �e�d���@��¡w�fc$��b��X���&R�
��f]�T��6�F�",oMG~�R��o�r>&�2�����X�`�ƶ��a#�f�MC@����,����I�3E)��sHfĉ>99��A0ok�����F��O�\E�W��4b!2�͞nOYMQ���0��&Y��V����t�T��?E-h���U���e��_	�Ƽ���8|�U���e��d9=���u��r��%t̓�@��܋�n焞RV��R/��kOT�>9�qY|j�yݏ��&����;q��b+}y[�k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�(@X~�H:����dܟz6O����p�(R\֎u�=7�7K�PO`�� \)��B/��Xy|�W�����z��3b��������U4����#=xeaZt�T����&�(���D� h�ҩΘ>9�qY|jT�3�7�*l״$(�>g��Ra])n#��;��L�ן���dܟz[���*1tSjv�[յ� \s�{��ҽ��q9+t�}!�`�(i3�����w�[�iK�D�b=:Xk��( fĉ>99��A0ok�����F��O�\E�W��4b!2�͞nOY�%t̓�@��0q�#�F��hd����!��R-hY�%Ͻ��Xy|�W
�Gr���%t̓�@��^́|�A���}o��Xy|�W,7��\���>��)����<�C,�#!+�+$�����z��l t�w�@�Ԁ����2|Q�-l�;�Kͽ<\��;��Cٯu�Xy|�W0/0`9N1s)l໶�,!�`�(i3!�`�(i3[:���[}�p[nۈ�d��-��!M�2*详p*�з=b~*��s��(R\֎u�{��b�b�*�eu�j�~ q��j�J^!�`�(i3!�`�(i3myC�0kc��g���Qrf�Va�ir��_~s�8	0X��f*��<<��lpЙMǿI?��g�F��6���xl�ݚ�Н�!�`�(i3{�d"���Uo�A��myC�0kc����Yzw�?0G.{T�2��8��Ս��%�r� ���!6�fcXy��q;_��y���D�f�.��!�`�(i3!�`�(i3!�`�(i3kǿ�E�Q�C��6�g�� ��-O$U���+���b�6��R#o�]�ʄ�;4�zu%��0q�#��m�jS����f���ø�Н�:���M��:�jOn}���ky!�`�(i3!�`�(i3!�`�(i3ݑ���&�d��ҟw���b�m��H3QAZ
0�1���~!�`�(i3!�`�(i3�r���h�0��X���&R���Gz�$	fcXy��q;ɕ�3_!k^���H> ��+�O�XÁT����d��-��!M�2*详p*�з=I�^$D����(R\֎u�{��b�b�*}2��L� q��j�J^!�`�(i3!�`�(i3��yb�	��q9���%�b~*��s�!*Ĭ����x��w����iK�D�b=`u0�F��aN��:��!�`�(i3!�`�(i33��0��|��sQ�G����)�
��V(MH��C��|���8!�|!��[](g���������lM�?L}�7�K��ȅ냇������iK�D�b=�u�w>G%�Ml
0j!�`�(i3!�`�(i3G!���e�w���ZxHk��k�z\b~*��s�02�okSbT��;�k2ќs\5 ���Uŗ�4�=+�Q��s�s�{��ҽ��d��-��!��KVט$����dܟz�X�R&cE���jVѭ@!�`�(i3!�`�(i3�N��W��fcXy��q;Pt��`���\�2��s���1�, ��-��h��Uo�A���x=��oQ2w���B}�����z��>!XM�#�yP��C��?�T'����0��d������h{���k���!�|D��J����1a�Hj���Z���$��U����e�����(�G�$�)�I�^$D��ү02�okSbT��;�k�K��x)�4��A妡��M/*�3�ܬ��H`�쮾�\�i\!�`�(i3!�`�(i3!�`�(i3p�@OM.Ir�嶬=���X���&R�l[�Ƶ���u��m�byBH�}�x&���Z����h{���k�XKH��Κ�d��-��!D���{X(���[0R=��7�Kc�P�z�1�rݓ�r���f1�.��N����k$ !�`�(i3!�`�(i3^	QW�Q!r|�;�Ojz�#�,t��B(㷾���E.t�