��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+��;:ӯJc��0"Y y��e��,w�*�iM{էA�w��%��
Z�ȰVo��������a043���v�ߊ���D�6�R65�<�!V����vV0��@�l�e��e^�Q_YYI�?��O�>���;�mOA�a{��A|�_s��#<�$f�n{ܦW��b�MQ�[����Гڞ7H=����(*��#�ԕ����8�s��(�>�&���Nx����7ғ�h-0�qE+. ��z�T��J8�����W��}��5g�?\��HS�j0 ��2�\�Qg��Z༂�A�z�DQv�DԐ%|�������vYx�-�F�h�Jҿfl:"�9�UH�6��<A����3�J��^�E�2�<�z���跫�?KacJ�mS$�����]�O0|,x�DJ#_����u*%s��(��b]@�5�$�Ӿ+&��rP{$c���7b�~l'�����V����ȹf�_4��W�[R����<�Ol�!�T�������\�鵍��27FM��=!BP�F���0��"~��\������k�_�^t��x�X�A���L޾)<n��o�jE;�\�zRl<��M_��gf"��":�,�D�ۗ���͝�ݢ+� �ځ�޷�|t�T�}_{Οw�4xy	��N�':�`��Yx��7��su.���b�w�#��m� ��Ϩ� ��������i��L݋e�c�Q=�^�s�3��qs51�xJ|�U�gJ+#�����.F �ف� ��vc��'!ϧ�]Hb%��.��P�28�}�����e��K����-�HRf�"��{�QL%|�@����6���+15���y(���p�:�B&�FH��T��?r=� n�Gu�׹������R��p��K*ⶳ�3���e_@��bEO�P���9|l`��_��L5��ݔ�1�]�]��5PK��ǽ�	
ǊyY��NT�X?��@p|Q}	Q�FAyh��z�A&�k�O�d�	�+cn�*m���TT��)��gu�p>�-���"=��EUl	�0�n|�}̽[uگ��B���OL-���3
c���F�Re�2Q��b��R�bC��uK�U��!D�_lOt�S�.q���_N�'o��n��J��������
,���:���v�D�GJŀ��#A�$KA\UU#p����gl�W
%�בUrO���&�����[Fl��Yb���< e��\&�E쇰+�5���� �b��;ws����H��ݾ�J����o��V�מ�o�;�,G2i�r���v�u[�F�x��h��4��)ɪ2�9
��=������u�(�|ɵ����Wt`���M9q���ꆃ3'C5?هr�w�
�D�[H7�8g�n-d�����@����8���j�c8k�
���!G��H��5CT��u��˰j��zXS��KS`�M����b��&��p<轐�р�E��e44z�3rD{,��Nk��KF:12��-�I�>���T�M��Pg����EP)Ycz�9L���Ixޣ+�3ަ�+�8���O֊cFx'��rq��͜����j3,��-f߿��7�^���������|�u&�h�'�1m�)��ˁt�I�I�M��ӯ�>�)0�Kw��_�Ll�>�UBg�l�]�^��*Bxw��q�IP�!��՜����t%�����*C15_Fy��+�k��M%pm�%�b_6�'�2C������y�7���=�2⭣����f����B�F���C(U����6g%<��M�S� ��D��(�&��P;EؕD{�5t¶ߖ���,�J�߭l<����>ՑvC<�+��l<��u���#�f��י�&g��_��E��g�'�����[����J#��
�#��k��Ж;����B��R�h����N�_缙ݜs-O�8x;�*(�0р�ko�A����~��v.����}�:6��Ǚ���缦�4��h6RW�J2>�Z'%9���E��2�ϩb�Y���g#�(<��cm�}���ye3���pezf���5�us��,��s<���n�(�ky�9;0&^s6з���5�.���s
�|
�s�HG�"��=s��:�%�#VR���:�xmj#� '�DE��I�:p	��2����IE����_�@�|�֎�>jgW�5��I��pJ'��.gSl��Pԃ��gof���d}ď	�Z�A,�H�$����,���Aq�-ڌ�z� z&�6�Se��-�A��Py��o��;��̰��x��(}�+(����'��j[Z��w3|��xT/q�,5Г�Oz������b(xr���(��[�#:�$޲g&�NVw{:Ǆ!�+�Г�`������1LЏ8��z�I�����j�3��3�	���n�O6{�x�B�{i��#�rr	����T�Z
TT:��%��J�3���J���e"K�@��8�.�:�B�?)8V�����+����T<~Y�\�(�����1�������MV�VIO�X�����!�9w�"�j"`�Sw�B���).RAPZ'~����41�sfp��i�%���Zjߴ�(q��)���k&!�;"���Ot�Hw��C���£���m���"_ B� (�kR��>`�������j��3$�X�ޏ%��jk,��K��#��Y��N�g��t��QL��1� �z�<�W63E�bq2*�(��f���9��t2�D��	\�N�A�zwֻ���ݓ#S���,T�}KiǬ������p��>}����uEG]4Џ���i&�cg�oɸ̴�I!�]8���e�E�� Y���d�8a0�;�I9��he+0b��GCә?*v��?��ް�k�ձ��y�� �ũ����c��L��mH"1������ 2B��GpN"��)L�U�@���[��K�qx�v ��`�	�w,6Uȱ��6��Q�l1�Q�|����ZU*���U?ƃ+�Y�
�Ǒ�<e�&�Z��JC��~�7���%�Rc9�S^l&�6�����n�!����}��.����wq,���}�5w�l1�`o֧��W�S���c;p��S.�o���#�=�;�f�f&���Ǚ2��4�ִ�ό�~����,�/������N�ׇ-V�F�m�{�Yw~>���t2�Z�@1�����x�佣����lnp�S㉶Z�4��A��7$�j���_l��
F��L�D�B���*��S���+M&(����4s"b��\�3zz����?�S�\6���#@Ƃ�b��'/�>�O��a�ex�/`�;��NZ�٪�o� ,�>Z�>R�J����h�k�7���	ᔲ�m�`�����[��@���I�`4��R��_�(���q�A_yre��f!*��lV5��D����4���U���;/iK��ƈ�t���6��A�c��LK�i��%�0u�����F���Fq��w�1O���zS� �p#���s��m��iA(e>��)�	6Y��ɹ�t��M�v�X��bL8�L�3���,[�3��"S�6W�az����#���@����b`�ۗ�!qk+&s��ci��e���e��q�q��0���}ݟ��
��=�d&x<�mˤ��pr#[D1tw�
Y�c�����|y��\�_Z�o[����ZG��ᜎUF~L�Y�h����46��� ��ԚC<o�ԍƁ���g`� �a�ט�X�� ��}�0���p�/C��~��|V�âlk�3C�x΂��N��Ϥ�v��Su1��ix5�Ž�m[1U�,��L�	�C�>zg������]	mF:������1���o;آ�Sq}ȵ�WGP��cg�!"�6�IO�Z8���/�Ȟ�cT�Z��]>$+��{#տN�������e��R�G�JZ�|�=�[I�uW�p}p�Io^,eaZ?��?^f�J�f
?�8ZP_�j�/�~Pا,�m k�H#�'�Um<�?��SA.tQw&���<Z���\İZ�0�=�x��j��V���8��E��q�h�DC(c	E�8g��q�l��(O�HqB��r#J1��4�'�Nr3>�X3���o�aL� |�X�ȋ���)2'��4�y��8��#A�&�6^���Hdڳ�<jx}9�Y��),��7���^C�I��9�W#'`�ߍ؄���TP';m���[��e��������Z#��̔��ܣ��}���88;:����Gٯ��