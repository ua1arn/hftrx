��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���Y�՝����@N�6�-�zi#�2yp3M�Li��U�~W�"X���ҿ��g�I��:5C�
"�s#'2��f
���
�Mg"�I����}+�a��!���㭍#h���-ɝ�P�:�B��24y�̮2�c$�u�̋��mƼ4��� ��>ٺ�a;%�:<Te�L33m\w���?9�8�����V�O�DTv1�S���V��ظ8��8J*b�<�T�W'AYnll(�aV��ʀ�	�m�Q�����������O��r
��@�A�BE�'��X����%Tj��"^�ٺ�h����7k�ݴ�M�0SV�*�@-t��Y�y���#X.߀���+G��#i{�%����9�f,��R�;� � {4�F����u��j���C��C�fO��r�q$����bK=MQjM�tP!��cv$t1��9>��r����(�,;G�>���tF Ќ�aC�����+ Q�W�~�LgcC:�R^�-�v��tm��0�ޡ5���J���=���ҒA�*��tef{�D�?I�	�x6$C��<F�[��O�k�5���>#��}[����7"��Q��2 ���N7���8O��Cs��~]���w\
��E�H2��I��ϋ��cf"�!9�K=�`3���_{������"��_��[�6&F5`�b�R�!&�>nz&����VL2�X��+S��~�%� ;��H�^>�u�ڴj��9��V�ܤ	Q@�^��o['����>��5�ބ�?z�D�� �v���g�W;�VaFy�.��0*�dԟ�T�~�R�r�c�O�]h���j�WVs�īή=�%�N���͛/]ƥWgZ��'ϑ�dAe-�TU���;節��ݧw��0^Z�~t��y�v+
 B�4���VօR[&m����{��i�p���w�H��a8M#��`<¤�VI"��.��܆�F���������N�ny���Dq�=�`�[��A��]��;�[���I&��.ܐ|�����7|��]^v0$ef� �͐�i(D7��q�17��+fg�����y�A�~b�WF>����]DV@�F�ē�卙R�i?�����m4u��s˯�����x`�C�۱9�$�g�1
7?&+�
ٛ4�c��('I�i�����_�X��+����L��X"C-�;�5�m~s<mv��_A�Ṿ�W���kP]�5�O�enU�>������0�'9�\�d"�l�j-:�QbL
ĨU����ݏ���iI�؃��u����K�r7���vI��h�m�3���U�@"(PVt|����H�����������c
��q��|ۆ�u�]G��\'�uʬ1a��HL&7�R�+`;3f3[��Ħ4G���@i�z߳��Zt���Pi��%�����/�������gV���*�V��,�l����T_!�O�7}!gn>S��ƀ�7H[{i��Ar.���b�o�P��Z�j� �S~,�i�"xՋeJ:���O�\��F���-�G%�e�� G��Z�m%�t�����o��]z���}.'}��\`8=���T�d����$9�0�Va>cu
��n���0��
��Cʹ�Z��D�.���zf#a)�u����vD�*�����FKP��u=ҍ,Kx2c�v�Q\�@
��Bv%ٲ�-�p�B�r� b�A"=��3~�ܭ��'�!��Rg����:2����GM�dt�E �w���^}w��r-p!��Ms֟�;r�����k��~�7o��f�.J�6�r�����'aDYMs��LpA_��������Fd9��
f�.�dlE�\��6��$�N����`�r�����R�)�ۗ�#�_;�R%��"�/��ŏ��[sE���1�W G�Q�B��ކ��}�S8_�	l#�-�X@H��,�&��V�u=m�IkƇ��U���P�֨��G��OB���|����˩e�>�v?���:ޱ͡�u���@�7�x�Iǎ�R�"���C�31d!JP3ҙ?�r�!b�{�*Y��c�m{<ڮ��Y