��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�Ck%���-Yڙ}VmCtT7=G�#�>�
پN��J��K�D8�ՠ�et�t�(�ӂ�&�;=����i���<��'Uj]��41��,N��ĩ���n�ӱ�(!��n���>������f��݇(��(n�ɍq8�~g������.�e{��J�қ�9V
����`Ћ$� ���7���ΑJ�(Bg����7�L�A�7�	�
>Ҟhչh<ti�����A�xm*��`c����j��?�)� ���rI���-K?YA:���qP杖N��ԭ���X��������A�s�I��;� <I�Mw��a�FγR����37iY�#�=�͢'���}WZ r�K��b�ml9������)�k���h��F�J��d)��-�]d��'h����Y��k�i�!��Sp1r���4����� �ӯ�{b'�镌�$p��ꬼ9�c�]�@�(A�������n_�� �G��B!\�u�wQ�����e� y�'nΟF~j��򜱈��F/(�	Q�3̯EA���H�>���^|����&R�GT�&Nb���D��뫧�¯&n�v�@,�5�]��.��A���V��+vբ���7H��O=�[��S4z&�#���9V�Q!J�C�a���Q��k1̝3+|x��y� �+�˾~X��}D�.��
��<x�������UR ��&O�oV��(���''�C�{��7ֳ��g��)�E�U�>f�r&d�,��ڟ:b�u��a5e�q�E��whx`�9x[�WU�net����؋u�CY��g�k(���*;'*;�P���� _,W�8��5�G�7�Dڭ;��vOD��5I�*�g
N�+֝���-η$ʰB�"��ʬ�D�s�Yva�uFÈ�=Ub}���G&}��J�����[i��������:�W5'��s�dE���+�nc���֛_��2���3J-�B�-?TK��.�ʯP LeJ�?�Pya[��K��)�I-劺Ps0MS(�j"M���ɒ�N#�����YLr������O�g��������\�>�~~7���̱
2@�ğ���$TV�P�F�A�G�ħ���Pp�&�/j: �"��O=����&$��}`�K��A���FQ0�RS?�(X�B-����n�`��������=5����LR(�h�������y�ON��HT�&�#�$����nO)N&�<.� �c1v���*j�,�'hИ���$&�1��h|.�µ��j;����oW?�L*��풩xo�Ϭ�%�o6��L��x��$�0H%!��sr4����^�;O����p��!�;�`|>�4M@�7�0��ӯ�î4=1�q����
����/� >m�
q����q��%M-���F<�.��a�9/�%d�Jo@s�1��]�zU�����T���p���]j;*O�n:�;͛������(�W��І錜�5=�S�D!����Q�A�"�q^�ZS0S� =��t�HT~�I�����hZ"@���Ь���K.�NT��T��9�u6�娣�<5=�~�(3�S��Qw���!m�-���NX���uH䇊��l�U�c�B�	�^���n�n6�F�)��Dݑ}���f��]���}x�nNK�n�C@ϗ���U��n_ȼ���b{��-���lK���X��4� 2�;�eM;#t��Z5�!@�,$��/��.I�By6���wpt~�~��C��M����Ƚȏ�s|Z�����4a.�[�;�91��$��܁C
[���~�"�Ǥ�``�����d�ɉp K�TL9��/��]�_i�����?����%w�.��vp�)���J򴍧��RL����YW�y5��{�ز���t�����ߑ �1�.8Ӌ���VIN�,)XנQN�3�t>K5.��pU���G�qö؉�
������^�*~�+�w�l����M���Uf�A�v��\���Ȯ�����\�@��k�ڃ�����$�t�����)i�Qf�$I8׶����OL�0�/�J.��=t���2l��bAWO�K�@���g��ߝ�1-	���)�=K�d�������$��Q3���>��B��=�Z��4^jD�#�q?a���vh�a[9`���q��s���e��[��-������!�� 3��7�HԜ�t��!X+� �Cv��L[�#vl �kߜX��I��n�4L��/�����H�u�.K{�C@��9K��3sH;���B�+�����u�ĉN�l���hu��*�[Jb[��j�����P>�4���=�@}�Z]�o��G�,P��R:��� �"i<P*��טu(`�h�!&j���gD�>.Q2�c #��M �g�wؿk&+����q��.y�<T����\��0�,����*_�:0ڪ��ۤ6¸�n<�磈��"$�^c/�]
�f��ðޛ�3��x��C&<��z9Wr�[��ȤN�@qi��Bx��N��T���k�:����.KǏ�E�B(&�	lo�U���mC�y�B����B�:���\QRh<:�.��KN�Q����/|k��p�ibKL$�Qm�턃KFu-p���wyv7ꍍB��q/5�TQ��T���j����/���o���چ�m.�i����9c�y�����r�d����6ϛ��Q+�`<a&�G���^T�ܛ$����T�E��O~u4����"��>R�*Zp�f��2�f����r��B����mƒ*��h,�� �����UHA֑m�$�vn�k�@�s����fpU�}yk�B�.�ٛQ@�'V�6�P�f	�@ƨB��Y���UCH!�4w��g�G�N8"v����7/���<�i�#���u��f<&��?�=����E*�\��!'Î�����gG�e�����U��#Qh*�u�'�q0�����S�o+<��~Sv�r� ��E�Q?{*s7��򮽂�'3�T�A&	.��N5�8���|82ք�\*U¦Z~��g�<[��"�.Yւ;����'go��mOPPb�?�
�d,u�)C�[������\Co
2VL6���X �����/��-�ai+F��Y�=k]�W�.jfW& N�V���8��'�wQ�r�
y�@k֚�S/Zx�\�󒟬�2�_C�g������d�+l��8�<;���4][�.�An&�C�(!��8�M�_�P~���Y�� �$���3���UV�A����9�K͙%����Ay��^'�@���?�͌�%��z�I�Z�� F(Wh� g*����l���ë7�C��9�BE��D>1��g��=-�,#���tɷ�{o�>�^���b2{w�0c�9G>�<���>�G��N�+Q�y�&GR���)d�XE/|�X;LH����1�/_�K{����p�a�\b*��@���n0� Q��j��@޿�z^�Ψ>��v�t|�~�ti��a�5����䄫QS|��ݟ�-`Jeɠ�[��J4�X�
F���?J �i>�m�a6���A}��+���&K�������x�� ��ꇻ�S�DU�@2���Ov�%�4�΍knH,Z#��>~��r��0I[_�e�62��:l�d��G����C�#������i�����q5��m@5m%,mf�k�޲���[g优��|[ܧ@0m�w��s0��眊Lǹ?e��"6^_b��g��)^�AD�ue�,�0�b?u�uܚh{]���*̢��8�Ң�c���I3qw�u�,�	V�C,��̴���-

ݡ�
��c�a����8 %������bom(� 5��#��c֨P�ҁ�W�أ�v�9��$g���i�EH���J���5�sv2R��
���o���N�����;�O86{�o�iY�� fH���>J���Ţ��
����9t3�A�	���2z����J�HL0�-�I�K2��������G�"������a,�#ް��x0ހ�RE�����py�2�d>t�m��c�
�}D�g��j��|� |�$!�gb-��8V��C49Yh���.r��GY$�yz��� ��0�H֚�p!?���U$�6�NoU���v3`�1 ������-���j�y�8M'����/��ɢ!ѹDT�jꩳ٣��
��=Dy٪�w4v��	sgO�[@��l�'��Ì�it�����ΡI\���5K��	���
��.�����p1��Fu7����1ܸ�}�1'��r>���֎=���OG����rj`H�*��ɬ�yy��Q;�ؠ�����-�� Ƿ
���J:�'I�o�E<���J?���J�u,x���(�~����G�;9J�b��J���$2>�toNt�oȋ��{� I�Jrl����i)�%��1�}�3�ec	^�9�1v�[ k'�F������ �g�ޟ��p=r�y�Gg�&��EW\��:+��ʡ�7�ʨ+Ù��3rz��5]/n�
��z�j	�Dŧx�۰�țŜWN�K-��R~?��J�:�e*b����3h.aߙ/3��|�{'f���A]���+���$���%g}c���<~�0�U���o���>�Y!Yn	f3�%챓
Ö ¢���iL
�=�B������1�s���2�i<'N�_���s������p��Т�
�ZK�W�1��Js=4�h�/=�c\ۯq{g��T߶.a���9������d#[E�X3�j�qsӷ��!o&����ž�л�3��F���lJv�_����0ؠ=w��Tŕ��p��J����8�u��������uwfX�޿��gh�6s,`�*�D��؍��mʢ\�X�.!��Ry�<��IX#�:iT�tp�������S����#ZTJ�֭0�k��Tуph{��Ư6X�J��W��j�N��х�d�ږ�U��dO�u�%��q���ףK�8_h�U�O��w�8}�:��yy�M��i�.����,/�!�С>(@�E���*��}��6�'��-�Q�ֲ�Y!=����~�������_ssCC��]*eҢ#G�Ķ/kZ��j8��n�7:"�C��l9uH�N��8�5��4L��)������7S�Y��_ܢ4S�jwu�j������x=����-5%65� ��#�ż�ණ��-�r���eA��[��cjT9\)�<p�2�2礪�Ld��ۻ��~�3��8�$.�3s�����-�����b�<ĥ	�8'{I��A s�u]J5X'r=�~w��[�f[�$1s�B�@����}�C���*�Az�r�Gã0�cM̜�\�=Q�
��a�H�e��P+���Iבz���\��څ��g�d�p� 7s��и�[1KWK�Y\^�[ۘ�pYFA�[U_���ae0���Rh��Ư���Î�*e.�S׃�vd;�I�hx­��M�qm��SVvS!��*[��t���$,�#n�(䜆���f[����v۰��(L�Gb
2R���E;r�Ǘ<���K32��N�kXF�z� N;`��B���V̯�י}�q%�`�&�׻�9b��D2�N! �o����mQ�>��;��k�	��� �#�� fM'�6�m��[U���v�����{_<�g�������K��|��1�t�id��F	����3O�ŻwIg�6���n�|6���\��EA	 �W�3'.��/�=y�u�t6�M�:�MSձ�	\���e��ğ����"&��iI,h�M�xrk��hb_99�H���"E�>A�uW`&��a匡�Q���x����v��d�Hb�I�6���P��:m]ˍG����D���e:�Ccd�����nBʫ�j�VvnV�p���.���U�KdS�� C����7LJh�QD���ep�{�RD�Cj{L��_��&}\�{�C��)p��Wyk���Of�6$�,r��ܒ���� �dC��$��r^&�yꅎ'���s*�1���r���Z�*��8}�O܀�N)���M�S�0:�,umz��xǄ�/�z�3f�<9�]I�s�����S!�����kg�~��ZP֖����/��=�ȗ9Q����KD��聐+�f ���F���޼|E݆�i�6�`t�D���R����CP�$?q�l�O�T-D�Wfu������G�� �ۗ���Ń-�<�;y����x_V/
s����k�R�]ڦٌ�Gs��<3B��wH���.�F��5�h����Mտ����$�r����&��=��/�Ѭa�u!�
"�Y�,Tr1I��)�A�/u7�k=�u3~�zJZ���d��W���nE��`�����O��+�ɛ���qFF����j��o}-�47D�-�kQ?�v�l����a���͆P*c�*���CVOu������!�0�2��ŸXa�)�;w�A����e	�����QgF�W��ne�w��s����s3���)<��Ɋl��@�.g[�{�\�BȯKΘ[��RR����p�� a�V	�H���g\qC���u˾M6?
��"CЁ�y'
&1� ��e��Cu�\��?��W�z����S��2���Zf~��7��i4"|?�(/J��n������8O����nʌi�5I���pD_|@fI3�Z_B�|�k�	�MMэt/80�ނ���F,�aи��{H@6ؽ(%5�u_�-���84D;&E�h�d@6���v������C>5�P���)�����h9�)6cꨯs?)���W>|�@��&�n�;��֡Ͼx�i.���g��D��-�dR���8�O	�22��2�L�K2�I���J�9#tC	����bQ��]W(@���_�R3�0P��L��fc�U�g�jm���t^l����, z�5��f���Di�EhsaK���02����}f�������WA�p�a����]�}7���J�Ɣۚ��p�H�+hp�!W�
��6�ԛ��iY�X뜷��Pp�6�!�u�	�:�MN�G_���L\Dr�Lɒ-���2FR�!�t���;�3���r2W�Dw�a��8H�yR�qZ{�0m�.�G���Z�T��#��W�̇X���ZN_4�JMƓ�[w���m��tpƵ����~+�v��D�j�6�O�ش�x�B��7~�/X{���g�7�H�(�y|�Χz�� �/~�_����_�:���e�D���B8�-��ؖ�|2'F����(v�گ�CŐ��3��~p�O���%�,�������TD�~5�P�m����s�崜@�B��R*�D��5x�����b�y}��F��M��g��Գ{��ܧ
U���G��9,��T����$���ֶ��!���Ѿ��9����a�F*?Ԉ]c\�n����ԛn��kj��Z���L9��ަ��{��:����p��h~�&vVuR�m��qǧ�6�Ϋ�Vޕ���/�mw��J9Ӿ}z{��n�<]��U=[)���! r����8�Ь�MXN3_��۹�^H �������%ڙ�~��}��Ŧ�7j17��GĖ�����<���U�.`ڇ�ZS;ɺ	��$�����zV���)�j�K�˻؜����jЈt5�l�J(D��'�˨2׸Ԇ�&b|q����ϥ���!);�vx&i�5ټ~veW����^A,�L��t��]�d�w�&�%�b��qg-���X�y|_�X��J
]�o��s]�5�>������X}�9��nl�6oG]4���^/��k��������i�|�;���ŵ+��/�{��Lϒ+K`H�/��N�u�oAa�"J7R.&��y��|��9_�>i�X`���mL���de[.~B��q�:����e���TRc�'.�d蕿�'�j/Ό��N/6`���&��}̱"�xVLk�?HM5��d�z̩�?Xg�zLevERb MRU��͔E'-�ߗ>�ʜ��jl�]�l\aW�|�!,��c��qS�%�}�c�}R� tWVJ���~-	����3P�@�KR�l4 ϹۖW�;V�G�I/`���N��%�%���BC�0'�b��QY�U��cN����F�%ʼ��d�&o"E��k̋K�m9�v���{�妙��(���$}��2�.5����{��\6��p��+��m���;a6�R�Jt�?�͆�+�s�j�O6fm�2[s��	N2,��1G�<6Wy.6i�v�c���1L쵘_���u��k�(��>�Q��ez5*]��"�]+����:���i�뵠a�����B^�ކa��Ԯ�݂�ˮ�ah{�]Ȟ�ԛ{��ύY=��O���I'��{D^&�õw'���0T;���<�=3�T-��%�eŽX�@l"� ږu���A�8yg�nN+K.��)m�x�&�d9�*�f�r�9.p��d `.�y�aC�M�?C��b`0��^̕ca�M�V�h����S�>Sl�G�@��m�l�� �D��!ʁG�l�D�\������;�/jَ�h�g�y�;�ܸ�H�}��0� ��##g��9���g�0X;�,���7 �t
�Sk����g@"�y��1Ѭd�ء\uU�N 2�W��ڝ�
�Nh��	��֚~�zNֳ�+���'��^A[/�+�|��?jU�h�A̰�����'/��=�R��#5�����]
A�0��Q�b��m%?J��u�?
���D�~3y���;�F���N���({xO�2?����'�V��$�Zv�D���W�	��4sxAeR[���CN_#�h\5[.��-S�v��Sدb��8=�ЎXǰ�`ϻ�R�zD�#��Y��?]�8rM�Z[N*S��s���'����$P�7Iu�U�xk�E�̼g�_��f	�y��F���e�!\0���\��&JA�$^�rZ^ȃ����(R6��H�i4��~��k�i�C�a9�&R�*Ҡ�֊]:h��<a�VYP���4+ߐ�h.5��C�I�[�T8 ��@o�%��V���d-�-	���~�r�b�=pN���c�����y�}���.#S=�-Ç<E�KT\���Њq��a������X�������P�Ky�qn��307/	J�g'쮇��u�#ȥ00lC����+%"��*I��$� ���7���1c�P�4afd�:G��9�Ī��U|qf[K�c�m4�;����^/�r��ܣ�f��������u����py�����DF?dt֋��?���'j��D����\`r��{=�f<׃�Mn 1	~������c�ݍz����՗�ƕ�<�� �e/��7�)�����0B��_��I#�9�L�m!��Xr!A�Ǫ1T��yf[�������&u�p\w�G�l��'����(^'G��*�̣�s�w��^�&$d��@�^i��w��+s�$�t�g�cf������]���f	t�A-��.�XѪ�q�H<w���+r��A�%��2c,ӿ�����Zeˣv,�N�,x�J.S �3rS�֖38|v�3�r��iQ���773��Gh|�!�x�fZ��&t���"��4�I:�m��K¼�����A͝<����d�
��
`^3��}�UѰ��_�Z+.�*鵀��RϾ�c���i��ش	�Ò���C��R�`�R
�c��ܯ�S�>V���Tb"}[�[��t��
+�:����;�����}/�2�������2��T��K�#2#�%$9q�%�G�P�T�j�+(�R�I[�f�s�PpoӓJ'�o�@*\�2�)BW��_l�D�7[�XG �G.^��G�CSn9������qXPJ��bU�ɬ�}�t���@��FFz<�"}��d����d��J�Cr��3O � !X��ˡ�`j��+�q��O�7QF�^a��*G��N�f��"(�:B󰚫��m�2y'�A4!^8��3�C��SZ��F��oAO'��Kȣ�μ4%�#�o��P�K���.ݵQS�i�	�>B��ܲ�ԞX����B���ʤ �2S,iTi&@a64��(�1p�!@�b04���7���]kh����C��d�������?����v��R�u�N�8��q�Rf��l������y/���dc�]΢������Խb�~�0_a J;?k.#L�����2��ߗ����3�����v�����dLv�?�D�#}c0��F��+�h�Ӯ��~בZ�/�eӔ4�?���8}Β�)�5�n�U��H��a�*<� �����$���,�<�X� U��X� �3}�3��:�1rK*'���7���9�x��  8.�z~BS�q��i���b�^<W=
�UJi}J��ރ'M��&�2�����n�[V�K��S��V�6~h�]9@^�H$�TF�!w�x��l��j����(ķ�WLgy!�r�����ߐ�c���y��0�ʏ���)خ���30����CApZ_���atʔ���H�y:o1�U+�0a�K7@������g-�(X�a;F��*��>��"�r���ۺ#j�ي���k*4m�e������_�q�"5��yXΎ�*�ո��J�}`M����S/��l�pi������~�Q�o�3]t��x$w��PR�K���(���կ�5���/���$�����+�3/�T�$���!���u8�ԯn���H�Ӌ�*<\,#����p!<4��I��V�	��g�ƻ���-�	����_�2�'��Ѣ�rz����ڪ���cϢ�JlWY_,`6e)מYV8����_�f��̲3�?O��5*oLD`?��{����~чm�1����R%��o�%�>TΈ��\��g#s>7R�->���7[)�4 h���Zp,WMNJ�
�2.�;������?;̥�5@��xy�\�p��~e��@{��fU����ep�[�Nf��	:j#c7�+L��A^*�ێ�s&�U����jT[�{�x��|N�������aAE�����ӥG9}����a�� �9&����jB6�Q/��\���k�)u�Bl&%��'ɬ�Nܑ2�RѲHL�n�j�Mo�	�>^�>�v~�[O�ۉ>Ov�W��8h4|�����U�rU��u��̻t���9R"�m�j����?�-�S���Bߧ�qV��X�R�5
��{���^a9�-�K��./�����<��о�7��֪����顽�g�#z'4b��� ��g�/E�l?)��Sz#��ª��΍#�hBʟ3�W(�~8��S�B0uD�������F䂎����J`��԰��qR����a�
O����\S{׳�f�J/�'b�q�px���"+e��i»�%z(���[S�4Z�"N�!��S�59���&]��8bZ0D�8�a��G��`��V����I��,v�Y�p��3�~-$�K���衟�io7�W1-Y	�Ɩv�c�o�K/z7]n�Xx0F4♡bn�
���dv#�#+r�}DR�%:���p��݊�؞G�T�-��\����PqH|�>�AN]�9pP&̋��u �H�e��E�r�6�v�����6bф�<����Z�y���~m��Ú
��:�%v���on���B{Aai	D 8z_��a�.����MZkw������x-)��3�z�\���ݤ�i���Z���?.N���I�yXKT}-FXh��}(�_�)EЧr�5�xH���f�}@�����lZ}�̙�0�8VѕA����T�՗��X2Z�ζe�X�j�Z�L��3���9�1U�-�4VV��ڂ��<1<���´1�K��J��	��>v�=�����?G��`�U��&`�*��sC��h17/�&����yi\�I�W� �c+�&n�'��8��ث(�����@Ξ��1�]��Yolq!���]���!��i�?L�Y`[&%�Pн�윅�}�^��jB.�7B�V��x��3<ڗ�$o/M�Yq�;a�k�N���魛
�w���R�����Y�o�ţ{������*()I�p2���-�񉏯O>��
u7��&����T4Kp��]����y:�+��*����4ӗX�y07�#c0�\�y��$�)bR!�S��}h�ݲI��r,hrJ2�����,�����W�.��{� � �XQ��;�3���'b�$� Do����ȖΣ�c�fM��A�b���fJ��w�"
*d�nS*�QW��H�^��~����T�z�z,��X��σ4����p�K<i�xh�i��[g�y�SH�S���z<�?V��n�L�.3h?��:a�Ώ\f�YM�V�[�+ �I̾�r�%���2�R�9/�G�����&�T�$g#9*t����Gx����'�h�ܐej�G��R_�F\�i�3~�U
/V�xa����嫉��8�`x��}4��Ii,_��Hg�z����4��˩,���6[�:����|S#�a��)Ш�LT��wH�����"�^���u���ً ��5�D?�K��o2ʝ�vju�f��L=������yr6	ݮ�h�����Y$� �[�*��n>T�U��=�'CTx�F�NyU���8Oa]��Mc�5��O�dUW������z�Љ����U�Aw���h��U��Q�ÿ�Ծ�2`��+K&%ՠ	�:��M��f#�K�L i�<��k�u3M�����x���H^�'�r\��@Fj�7��U��\�b�	WM���0�������W�(��Cq1�Z~Ɓ�t`	���`x�E������A�����߇��E	��!��ix����$@���2�3D�_����G?������CѺ{�at�W�M�<�|.�N,�W�*��s�+�9��T@\�3�nx�*��o�Q�����ҁН�,��p��26������'��?�����d��27�;�������>���F�d;����S�1����Z�.<�0�cr�p�b����o7®v�:	���)=��:$j)���Kz9��*y�3����S#��%7t���ʤ����/4_����I���e�ƍ5a���`���vM,��~�ѝ:���p��Y�I92��� �]��d�%4��ߝC��y��Z}�u�Y-�s�E�p�`=,v�NRؖH�e�j]/�	F�,aO��Ȅ�>�[��#G�%�J��/z���[z�o+tu�ث<�I�!����),�4啾���p�,r��/����u��F�b]���I�^�(���=.�[�CWе�T�?��s�Y��.ƲK-N����±��yQ@��`�';tO�K��y���~Gޚ��͝�:�,6�����=	q�ۃ9°`��has��[��m"�H��%~ ~��; \�^�����8Wu���R֔��0:t\�	NK�a�ym/[%x��f�鲙������@S��{`gQ(Q/b�!8��n�� d���038���yFG(I�[L�ܔ���Z���q��a�%���͚oJ ��Ly�َ�������Sa�&���"��l��V�./�E�|'�-4��b�����b@�D��R�jm/>�P��IT�'�Eg�������s�`�~m�Ҋ[���������З���P�`�?�!�Z��.����ƞ>��K�K,�����j֋-;L����v�2�ԩTZ�����mŀ*���*�H�e|=$�J�5N�a  /|�����u*P+؄g���c�HaFf8�6����-�o.-yU�.R� *{L�ÅR�#����e������F[�	�z�",�Tl���j,"�����b"tz�I�@f���RTM�>�����P�"T�2% T2�v/L@�V�(���E-����lW3ő�|�?��tH�|�Վ �_��{�Ʒ�n����"8�G ����@��qף[f�b}��@T��tS��܋,�$�{R������<��v���?��D�"�C�xߖ��3��kW��0w�H�B��5�d�6�
�Uy̬�m�8Aٞ���"���$���e%^�Q)ڟ��.,ťǉ�>w-;h�{�8�X;KP�9��׹�7I����a��:'�G'�� �ߣ�9��9���QAm��Ϫ���V�֫����(P�I�U"��
l���,M�������VY��`�}:�պ?��O��3y`���l*�P�$S.)��φ �֙�!���S
�L'�N���nvNۮ����_9X��rV` V���޳.��͎�l��d�d��Iզ��|���)����^������D<U(,��P{�e���q�eԖCPr�ݨ�1$!�������"�£Ӈ{KD)S`�÷w\����uۖj��0m���I� ��s��4G��-���<���uʥ���ϧ�0��n2�w�S�d٦�[]A��o��`���#�F1�XV�|� ����#�n3���-�a���e,�NǃXI���~��*�*5a��Oy�G�6�#�/��g����$���)?��p'�^-��8`kT�UO�g��w�+�l�`�j )!� 
��4��mZ�5��)8�v\�-#? ������>j����JFAރ�o��q¨�v��l�����}�ʄ��x�D��Y݅�' ���qݧ���2���=�TGF��ՑxE֩x�.s`�"��:���W��tL ��f���z�^{U��|9p�v�a�9ܒ��|+*�}�+����3w�;� ���"�v��C�>y�qr%�|��T��3wQ���������n��<�BR�e�-�W��|]�Y�O��-�e�6����șzZ�m�̈�'=�$�����GB������(�|Rt��Ȏũ�N�G�K�I��Y���_F}H?����[7��8�6��ڭ؉�IpL��t�>,��p����!�j��#+�:�e��,���Z�*���/�gI�9�9�(�z�So��)���}+���Q]-��y��pW*M�ӡ=������մ��۹�#U�?�0ǝR�1s�.�&e�g������L����(����o���U'����|`k��|lS:�~�{�ul�[I��!6�?U���_+Nx��q�[�5먟`�j<�$	��gx�[�H;�ǙXj�߻�����y���!��yc�~(���O !���X�W�f�Ce��wl�ƋCrG���Q^<�4f�.�<��i���S3ݫ�%���f�cD������	vC���&s:�p��f�RI�٬6���`6�HIo�|�)��S�~�K)��O���󫢑�7�Oc�j��ID.�B����,����*s�Y�\�4zSz��*5~�L�?|Z�uVp�l5� �h��g��F�+ �&�)�^���E�^��
{��+{='N�n���9��4��L�9Wj�zۊ� ���)0������+1����}d�4ȇ�鹗��ai�Ɲ�wC�C�y��G�iHe��_�&���%ٗ�Jt�7�^�.����%G�}Hɔ�k��x�͏��Ln��߱����� �ڻ�����z�S�칀�q=��Y�af��z�Z��'�z
��@V ���n�����P(6@=jQR���|�~�Xn�ґ�A�uc��;"��;�֕�Н��|z�{-�F��b��W��QG�k�'	:y;w�u�,7�vES��c�}Dp~�r���C^T��>�{Sy��ݧ�&�/�G�|�3���{R:^��&琘L�m���e��p���`r�R��W0b�^�ݏ��p-�zW� L����F?�[Xn2)�6�Z��/'��kqý6�x"b��]�SL�e�\2m�������P"wv�_�2}�+O���TgV0�eSƭ�Nb+I&^O6�P�6��%cq���qG���&$���*ĝY����[W�K������)���� 9����)�Qnq��@�J���d&���$ٵu��44�6�ORCBD_�<,�TZ�!�<��5o_L��d�@��މ�Ԗd��Uy�d���Vg1�1�}z��S|��6��_˒�_Ɏ��љ���|�r��H9�W.�U4�(��Ƣ(�q�x�f��m��7��F���#E	�i�)�& � K�����!&k_ĬbbG�~�Vz
��L�z�
b��/E�y���eU����,r�s���)���>?4 �(׌&�K�A����+<�L���rܮH�����.�k�.R*w��m������ R��&e|8��*��`N�]wnj����Y�3�,$ \�2߶��a�����9N����!���q��S�e>c������?��@�ȳ��;��?Î2^A�YM���nD1�2�U�o6KF�
\�4Г�&ע�I-,�#��`��d�$mw*h͐�{����=���Oċ|pm=|��T�d�����w�ɅR_���B�ysd@�a��`��E���z�T���ܤ���@��2��N�Ҍb���;�wf| ��je��<~�[s�Cb�Wx҄\�
�n�\z��^9��������������jH����tɄ�Ȱ�s�K���A	m�<��@��h��{�骭z�<g��*�c㩳x;��d�F@0N��L`ԃ�r�@֠RQ5�@g�L#���͇s��"���(�ĩbF�t{���*>N�ϋ��a�9�|���n3%�)�4�k��_�l}�5s��l�ғC+Pj����j�Q6��,� �o\��=Kk1���J�o=9��۱��\��Z>����5i��#��7t2�b��H�f$X�$JV-n'��"���R�yvz_.H$f�K��C�L�K�<��[?���ߨ��&�j�7걨䦅" .mQ���y}�����=��bQ�Ն�D�1h��#�D,2����f0�`ߦ��]̩�-Ko��������f1nGD����)��ɛSu��'��j�-�
9<d䬕��,����@�$|�9=M_�����9V0���薅��N�̠��Y=�ሠ�����h�y��b�aQ�l�w�Ά�,�K�p .=C��e8����+_xu%D�-��{]M��j��`�>l,�F��}L��2wb�i/��}���!h�zM(_����m�����nc��
b6>c����`�gl���l�P��+r�(|���~�>��t�]vG������i�/b���G)ګ~�����=��������8�5M�9��Б�/�2�_��7���>_BS��_�Dp�>����V���a�u�	�ߡiUg���X���-dߕ]/�J>Q�q� vz- ���~��#2o~*��>*�2a�"��zP�%���)vR�dG�r��>!I�ތ:g�y�ըf�HfQLNqZA�cB�eh���O��{^2�[:]+B��9��j����$'͋�؟o�1�q+�,�$���
&�(3z�X�J�ã�'Рp�Q8�������M?��,�@9�iR+)�L�M�O'p&�J=-��BaB����cU)Т^��3�u���&��ud�ЦQko�?��~��7I˓Ҋ[��u"5�^��ެΥś�ϵގ��u�diO[��?E-�����y��o�E����o�~�[jo���(1�jE�TP��}躷i�YVs���3��ZYb��WZex����A/�pi�����g$��K��0Y��x�I\iEF)�b�⏄Ԉyg`�9X�c�'�}C�bj�_��M�1�	�NE�,ɑj��L��K��\�~� �Q|�8@r�!���?~о��Ł6���
�~?��r�)�{�Iw�([٬��ۺ�ˀ�,�ڴ,�'��Ft!*����5mv��F�*=$�>�"��z���'�:*6uBE�����	�Z�jy��@|���_���U,�+8s��o'��,i��p�C� ���Ӕ�T(����σ����3�r4�G}\�g�iJ���&(�l8p������Q�R�̡�߮��m�7�R0Ȝ�w�&|$�uMn8��2�d�isv"w�����c��G�T@E�]3=1� e�(��}Ku����T�tg{��*�������
����yuI���O,S��.�,�M�u��I� -c��6�E�E����i�I�)�A�n�+�+c dV��[�D�V���"N���!D>���W��؍$��t������y��v�y���Ut�ݤ�e4;����i+��E�ٔ�2�j���=Qi�{տ�;pL���'bc����y��8x#��l;�g����
���0��oE�fouj�oz��3I}^���>�N0-��ݯr�8r���etM�DT���7SH`��c}\�B�B��@3�'�=H!��n!��V����u�6�5�Ui!�Sޖ8_�ԉ�2ۗ}�㙂P��y���hrnB$π2�0$���>|���Xt�(�{v�l��*vZ�H~�a����� ��l��3$�2(L	!�y��qc�R���Z|�+R�J�u���������b�}@5�8�-�(@9�$h�{�'���k��3��B�ck��fDt�����HM�h�l��w+t����r�-�59��� J��6lI���!����c����(��^�>4vuR�7%����| �������Dۊ����aN��6���k�Z�^�S��ɺ�)�kp�L�-dUu��ugo���h�� ��SF����4�5C�D��ڞ|n�	y DG�ٸ^f��kk93{�fR2��n��� v�f���W���@��'����ݙ!T��O�����{��a7��[����#Ր�9ʁ��?4�3h�u���NP�",co�B�8.C�}��;8^O��Sk҈�� ��������]C��@��+�gtո�9�²��Vm�{l4kC��T�h� S�߰�������& S�����7'��3��oj�~���7|�-Ow�O��+��/����������ZT<r�Y�o8���P�&U�h`-�y��N�v/��� ��-���p�4�d߀�:`=��D(G#�P�����4��h;4,7ho��W\ނ�x<�O����B@���n+j��3�`��H K���@ԕ7b���ւ����k���,AA�h8���j�F)�R��s[����]�Ӊm�5���{v�M=�U�8��e@����{�~TP�����߾
~W���n�Z�?�՛� ��t�����q˦f
�'��}�$��.�⢢�D���u\<M���x�n�j�*������+��~o��э<���z�IM������`� �`�ƊSz��T�Y���Xr�
s+R�B�o0a)Ks#A��R�1MR;Bۗl���AġQ�4!Pek�ݬ�}��e�%��M!�����2̐ҭq��5��h�"4@�;�n�Cu��ii<��́p5�*T,���5�*T	�P��������L�53H�f�4TD μ~<3�x�`lo�h.��y���l�`����z%�oXޟ��h:F���3��xS;���݌NT$`�B�͖W�K�����CHۃ`
W%��'�j �}ჰ�bj��Nï��!x+���B!6�'?����tLq`4çv���$�Q�\FFr�?�HEu/�E,�n��_W �P��I���� [;`����f���`�C#�-w�oSvY�^�ʹ��*�LLdd�5!��c�e�E��}���j����Z�_���n�o���������hP�=mN�ء�vSKƱ���ln�.(4�,��������5?VWj�]���Δ���)�Gt����	7��k�Kl��*��R�Ǎ�:�` �'���S��ۙ�v�Dq���ݼ�/��Ez�V�39��ʞ�9�,_����Zg�{Ձ�nI3���W� v����hx(9��	5]�P���(���ଏ9����%���̓�`�r%����C�%忦F�[��x@B�4��-�V�7�[�1EX����۷$�lF
s��15�ͫg�Ja5�M��DQ�u���WU�u�Z�s����t���S���=�'2-+'r�'�H�>���0gK�bŔ�g�-Խ�F���!���&8K�!g��M:��:|(�g�\�f�R_FJφf�u�W/���ou#L�F|�d���y�;N����f*\:I�h�����͈�;�U!"�C����|}���I�i�r�f_ߚ��)+�)��į�KIz��m@7"0�Kw^��<�qG�Ч��x��PxvN��#k8<wx�+ 2�:�Q���N�oBDݩ%+]@�B����0gAIh]{�4b��5�+��z]�۩A��̼k-ܲX^>J��0���WoG^ƜLD�%u�|������HbW"�Q�ʘ�u�9��}�IR"��m���Z�^��]���\���)n}k�X�-��U,!���D]�^c������ʻ�FzvL�.C�B�m!�����=�"�*��NQ�Ǳ.I��͋6g��j�I���X��bQ({��X��îjw��yԯf\:�S���a���;��?������B��ď��KqW����|���V�7؆V�2/�vb��M�,�b&�3��x�j�P�ڄ!EWV_�������>E{�*rvOh�3��྽�Hs�DӏK�dm��(bx2���_�=.��"�,���r��>�UJ�II#9/�֡ԓ�j��8����D��!�eU���� �k̢���w_k�r�/`�m��	r2,!K�#�������A/�W 6�p�a��fx� v�=h�2�&n=R��+�	N>�8j_	�]��4�*�����w���CJ��3ga=��9D�х�Rp��;�e��P`�k��'���w�� �hR`¹Ҙ��S����ؑ��u�+�V�~��-
����b�s�+�px�DpW-D(#�ݑ-Ǘ���ZE[����}[��+��̀�ܭ�V}����N��1%��?�m�g�X�vF�k���a���&eHEfE�N��H)�pr>��7Jb��M��?,����o�M�%�<M7�i��V���K؆�Q��t���B�
Q�2y>\� WF����t��;�H��C�Y�����R��I�B�DE;�L���US���6�:|���Z���TPr���}���X?������?�z=N��������.qGI-P�������r��b]x�Q�e"�V\��=�Kh���A]����Ղ�����Y5���DD���1����Y}�y@ȿ���	 Z;�� ��E�VGՏ��Z϶���[V�`��B��'�q|܁���9����f*s�(i�)g���I	ވ�xG��v��Dk�W��UH.�������P`�"�Ja>ϥD���c��++L	α��f�����^j Ӄ�����'�мB���K���ͮ�N��h��Ulgop�����?]�"�E�KV�u��^�@o��h��Z�P`r0�HyVk?��,>�ݎ�̈́r[��VO�Q &,�a3�w�ǧ�W���EF�̘�|J2�n���P�W�� ������y5���i�?j����س��9���E��R�5��ȇ�0X��. ���X���y��������M���bXK�m��b��gw�\1�J�^ `��}��PuW�$>g�}�����wR�+�aq����¼�/�~	�rsG7��$R��vʱ�kah��;|[��@�:�L]Vi���r{U-�����=��
r�����T��e!�EAL^n�����~q}��s@]�X�!�;�Z�&��AZ�Նq"t �V1(�ˀ�H�.���h��NB%v6.\����[�|�5�b.i�������CU&"^J:S"��d��X΂���� J��xi�Y�#�����V���Ϧ%n8���5`p����Eg+r/B)<V,?3_����'R�����R��x�y��]I4ϮާU
�5�$8u
CI(i���	S����㺟���ݔ�:Ҵ��O��[�T,���z�v�4�g48\ڗ�ru�Q~�������`7�J1kӏ�gz��K��sܘ�nz���y��>�Bp��� �-���,�,-��<֛�}~n�fJ����QZ��������"Ǆ��[�d���2N�oa=O.g
�
�)�fҢ3'+��Gƕd�p1�ݗ�	.ݐ6Xp������Ӏ��ܔ���)kt��p�;��r#��Y�����Ϋ%dlk"+O�exxXt�Ӫ�ݩ���<?@nt��ӛ:�P���oQ�+���h۔lSe���-/��(��g�[��YTjxjf�,������t�(Q07;������Mui��&��w�5�[�僾���]|N�W����FC1����a0��bV"ёS_>Θ�����.}��d?<����s�J���=�����.�,��[�FAA�dȏ�r��	N1B٢B�U�X�L\�4�29]�I|����-3@�Ձ�vohgP^�נ��Ck��E4✡xE9RBć�^�ݵg�����W)����η�^�}��x��$��M��$�3�V}B���>��P�*�Z7�Zd~|R�G������!f9fiF�;y�{�8�<�	���3�G~n��J�1T|�ΉrR1���V�_�n�8<�����l�z�p϶��*�DM��T����d����2I�C>�:o��o<M��l����9?ɱҋ��Im�Oا�d@"f4��3��C��G^��2J����%�uaO�X�T�H\��eo���,]�6tl[�Lr/��G�AŵYDD��/��v�'�� ������쒊��6���+|]<{��2<)�� ��В���;����1�(2�+K+L�j9����t�*�-/�a�>��bp��ϔD�7����+RŲ�� Z����D����4�S��K��sװ�FV|0��V���
O�h=�d���ϲ	Yo��{��z�)&�ݺw��)�<Bn�~E8@��r���Xi_�!s1
�#��O� $U�G�D�S�;�՚, ��T� � $X	�z�8.+�&��<�J<bq��`=Nf�N��m���s����5w��j ʗξ�V�L��I��vR�l�Wg�aɁ�P?�}�7v�Ƙa�k���5��Z�!�&s"ƓS{u!��uF���aq������P���N6�\&Oe���:��.���"��4��v�b��{�P��>'�x�|�iN��b��������1�EH��#W]��o��l�O�GC�j��_� �"#v����jo��S�Z_˻/�ZF�kDR����ῩY��۩�}�C�Љ�bj|��|�|  �X^�2E�I>O�'��*������.##g�D]bi1:!x�!'vQlC`@mV���us����r�X�#��6���v�$��Wq����&�X�}��5~#�T.}�V(<V�� +l�"6a>qGȟ�*�Q�֓Wc ���M��n/����a����c����*	eO5����jDD��=i�3b���<�-)����1&�i�u�.�U�������=_v�G�C/l�m*筤�����u��b��5*�猿���f��4$Ǻ~�2��f*���
Hj�ܴ��5����G,�k5~9)��o���\����^D�������7/�}��ԴC�}���~�<��Ln$k��P�l7z�,�?Prd����?�#b�~��їY��Չ���43�;�%�L������eZ(M��;��C�T��_�b���r��	�[�2���1��?n;�Y�+FE�Gy��qV�u�1������E��l'�0x�ij��OQ�D1XQ��N�N��L�z3�?(�
?ݢ��`�P��6��ƿ����?�E����5��t�ĖDj58��ڄ��3U��߶�h3㵠�jbN9�A�#*��׀U#Ô�Q�ۿ��.�hV�R�Š����ȆKdrk���VЂPm��ۂ
������T�G��|�,L*vb	/��_��O���ˡ�AȭI��?�u���5���}������KK�]+�&V���mY��!_�I~��?���}TE��Qh�qg������ƹL��?SY˭�B�Pu�.�a���hm�%\ �4��4��F<���h*���4<2J��,�۠j�mc,�I�ykY���A1���+�������:\|}�#��O��yQ�<܌��Jw�1q^`rv��Sz�����@s����J��-��%>t�N �s��f;�
0�ǆ��,Q��o�����"����{���>5
Ɯ!�3�z#R�����[j�*�P>m{>�g�	�H�8%�h|��n�<��/��\�`���vT+�јV��+��I���������t���l��w2�(y+��] �g �+#
�D	���C7tciN�|;����!���Y�ct����V� ���DQ�óqg��*�S�!�`Y���+�^���J�p�Lh��r.�
u�y��&��	�gO�n��������������z��y�n$�J��ϝ�ӳ�-y���j��u7�_��;Tu�?� ��<�~�ր��Cʐ!
�KI��'��ϓ"���/<2��~Lq�$�8dILC^2�>��"k�7��l�uQ0�Mo�������)��3a��?�#� ?`�,U���k-u����?�L����P��3Y���O̙4��?�P٫ٵ��n��Ş/�"	w9=��q
��y[�/����$k���<�,������6�t�7|�Uwc ֍O|f��2�hL���c"�;�$m�<��VtT��ݴ�����1R굥~�ݟ�0�����<�Ze5���su�U]]}S�b�8��><�U�:�mnD�kz	`Ap?�f8[�SS��WS�gE%Tn���Pz�ǣZFGU�8t��H��ֆ5@�6!���2��e�<޺	�3����b�ZF�9[U��� o�X����YS �CW�,�%��k�I���!C��ܓh�b�]��#E3��Vf�x��5nrO���
�]+8_ÞVi�}���Ks�AI�����^�wT
(h)��5��N��bڭt�����غ�S�����'�	���ta�X�ٕ&�dy����yjR�I�<Ή��.3G��F�<�\xe����X���8Nt����{\'L�ض�jZ�M����T̘��If����G#T(���x<P����]G�#��|>�Pq �vy���4��F��2��R�.p����ZQ��2eTenf�(~>�i��E8�آ�A�a,��	MMĝzڔ��r�f>��'���Wٱ�)D�Y�J��އ��'�']Fyzr��䍘t+��=���1�*M�<( ���6�*q��"��|���Y�U�S�eOUs�1�ghJ�d�����b%B8<�j�zc�S��8y�TB�VT(�T�A]M�nЉOe���.i&"
L����Y����D��I3wG���-A�Hl�67�	�dѰ������J�<4�Vp�h�/��B��
a�e�F��zA �G�c�E��k��������a�!9uK�=ҥ�7^tzƞ�4�*-�(f�+�D�F4!�����io2o�M� M�Љ�ܵ���9�����;�,�?�IH}>a�Ѕ(;Kj����%��L� �ے_�M�+���RI^"p�Xj�JZ������\7K&ۈ��K��lv����i��7C%%��lm�f�ƈ���U�"GA�rq�l��9��M��xϧ�m�{2<��Y���R�y��#�t�>�<���!J��X�&H����c]{g�Z�#�4��i�=���6J���-�ҸWm���re9̤�=�&z�uu�YE�ǌ��Q)����V�� ��2�!S�Y�Z~���.[,vw�
��183�����?�P9��,I��mX\s}cг�L
&��'�G	c��D�����w�Y��yG:�X�U���(A�>|��X�x?\��
@G �!��M
�o'\��ތ'��sH�nd�G�Zv����v
���)��Q^ ,�'�ү�t\`���w��4~Ȧ��U� ��$m�sf>�s�H����oR�3��=UW�`4�eEaz��(+f���Nd"��6��~c?��a� ���� 2������@�aV$���w�\�釖����4�?��S��|Ѻ����T�,*��i4�l֚����%c���ϥ���v�2�f��>f �A�Ü�I�nr=�ߔ��usV��n��g_�e+@'��{��\�X�%}^Ƕ��΅�q���Eu���ޒ�wv�e,_@Q��@���8ڒ��l:�ń>�����[r��K3��{�p2͋x�z�l�G,f��{�����E��6J|k+ㇹ(��j)bl��N~�u�jہ��\>P���{�m��oQ�b���(�d��:@��X�5����r�=!1��0��ԡ����p]�e���e�βX/z�ƞ�Mq~�&�!b��`�u���	�L����ZԳs?���|w~j5�f�X�u[�P�[��������ͣI��I��ϝ�[3�����"�9HZ~��s^��W���p�n�@K��.�����rF�h|Fr=b>�k�0�R�>&�$����nbB��!hyy�Y��֏I��at��7�a5#���a��h\{���f��1T�my���!'�(ùO2�=�����u�R��	�5��:���x %��Qp�z�d��H�c��N5� ��z��:�jRҘ_�h���a�����y�H���R�ڷ��X��2�r��RK��;󻙥l��(�*'T��$ �nA�m�i��\��,)�=��cH_B$7���6u��q�ȡ��f}?�YQQ���}���1�J���Om@pZ���ޝ!�xG�V��R�)���:���"����W��ClҊ�J��wbVZfg����կ2v��կq/a\��C�L��]�ga7�DE����<�4�/N�mF�O���}��ڒ<�������̠�qPs?��n@�����(�]����X��C���C�����^�MLi���wF���rCٟd�u���V�I�K��YMbԤ��$j�+{0g�
3���}��.T䦟:�Rk�v��PI��6�e����m:!"�0o�)�U�_(�8�����GroA�|`'xa4����%Ǿh�4F�p'-����G��_z��i0:�*<L�Y�h�5�y����I���1��U�n��_P�ʣ}�Lbj�~kD�4�߽)d�U3�� ����0hl�<�D���(k�a�bԞ�����3j�?1<\�©o ���t{�h��J�����%��f# ��`�ⷽMiZ-�����e/�j��9���	��2��cCE��N��V����*�o*W���'(��t�W��Ļi�s��u���&�{9�-k`!"C�)ON�H��σ6��ň�v��@|U�C��IR���7��"��5h4��;�"�R����8"���7te��؆��Ǆ$<fp&�
7%M�qJ~Mxt���c��a�������;���"�R|F��T�p��s~����:���{b���Vc��Q羫pn���9���S�@]xN��$Z1����CxRG�ʹ������.���D��	n��[*��W	�Id��#b�e�ðJ����P�������>M2HR�ӦZ��,�J��xܑ4^�R��Ĝ]46�Gj�1}}�����8z�Ȯ�w�3�����1ş��E�!`^�����L�� ��l�$v�J� ��=��JЪ,�g�_��|j_<K�Qo�$K�]�:�۰�E�x\Fx���o��@������ȣ;U���jL��h�ڿ������h�����#I��n"��q$�=����}Y{=����p���z!�D����S!�;3+&�/k���F�Q�j^�w�;鎯	2����#�ށyN���@S�f�lN��1�o�{�����L@���.��mp�����,r�B���0ŭzV�q���x\��lպc���Eţ2`�<�=� &�U���ИV��"6��'ߠ��SݹO�� t���K&F��kR��UGlp���IN˽J��a�����Ok@Ͻn�[ʑ^����R_f|ߣc�|�ޯ��7��w]24�}��	�q�֌>h�AGں�$��]Uu[���p/T�
��V�Y �IY��5'��'�;�w�IWx0�G��%q(s��Ye�Q�����|e�[��'7�십׌���9�����q3M2�C����º�)r߿�*�b����7�ֳ�'Hؑ@�RJ���A
}��6�3�ɓK�k}�G�x-he{Q�〄�`���M���z��ә������"H�g�QΝ	�+�$(W�(F]�m�A,���D�iKGc�j	�5�t��E�ު+��Z�㳮�r=hi��`N�W	�*�?V1i�r�>�����1D� �0�e��z�Soڬ�L9��S��-׷F"TkU);mB{�Յ�=��h�^�9`gV���.���k�z,[�z��i���7Ur��kW7�YcЩ�׿���Oe�RQz+��mr(#�G@�h�a.��@�WjG߇�� �4��q�4	b��ו��h��d�;��d� 7}� �����_�?��\|k�;��"Ѭ_�))���]��,F���L��,;�����'X�<XӚ�����{���-��LQY��SAz0���ai�ۈ�d4�]��w���m�BͷKx���%e&����9�x�R5��|��2���:�L���� |+o��d�4l�� >t%"���4Q���,MR�0;�cW2�lyČ��V'�^��N������Q�bߚG5fc��|-t�r���U�@F��m4��5.�)Ht�`�|E���Ч�[v���?0;Dae�R$��K.��}q{��[Cc&��e�n�����>n��N�+�e������mx;�D������C"XZf����S�\�>��3���� �p�z�)+�d���@��bi�:��9�γI����[�!6X�$b<��F�#@OU��4>'W�"X�al��M��e_ޛ�t��3Kǧ��$�y�S�ߩ�/��{ܳ;K����h!�%���b����NBZx3S���G0y��&�fȬ6W��b���h�S�)��+R �9pg�&P��ޖ���eUq�Hk'�g���$tkn�ea��w^LE��Wb�{��qx/�MŘ_�4�(�k1;n����?tT<lm�d�u�j�
i��|�!1�Ɯ�T��������9Ov�7���ۈ��c�=(\�X����� ��R�}Z3�-�C�h�g's~a��d�t�v����,L��2�N�Ek.	���ni��E�����Oy�4R�������cYW���)�??6�˜�`�y J!�uE�O�����7|�^�Y��_���+d�x�,#���cˇ@��B��"4��y���>�`i�2�O8�������I�H�_L�rY喊Sc��y�{_ �!#'�]Q��W�5H|�c����YͶ�v��X���^�X';�+���"rbt����u�G��,"\Y|0���$�$p�H����va�r�3lXߣ�G�K�Xg�(��Gr��WN}!u2iw&�3Pnu�u���ZM�SfGi΃\�J��?�W�T�@�Tk&�S�NF�8?���Oo���":$j?�p`��,�R,)����S��Z3Z�U*+�\..޲�˵��5�ny用(	�}J��i�e�n�Wk1���9��m������ȦX�-q꘍摅E��ҧ��!]
3������Ȫ�V��g�ș�%�I���%$A.,���13�p��lZp�Cd<�P�$��!��a��O��^��긚q�c����r?��=���Q�c� �e �D�z�β���)���ul��Ӈ�T����W���[5��Q�άf�H9]�l��ym��\ވ��b��I{�Ki��-��r�_ٰ�}Qo��=q�sj���h���+��#O���K2�������E�}8^k�Z��И�c��տ�2���x"�n���/����_ ]Gc�$Ժ�j�ncy a�R��ݻ�Æ�Z���v7O�u��֭|k)�|�#zp	�� ��F\����
l8	a�nH�:����-������9�T�/�ظ-���E1٦gh{�M��(���6J*�>�<�%RUfn��1G����;H�i&�*������9%����l_c�8�"_O���]{���#�����b�&�a�r�tj�E@ф޼Oˋ[��*�r�R.d�1��[!��(2��FK�2�}\zn�K��i= �P�]�^�i:�X�Z㑵�\�4`��)i�$"���6�E/���eED�M�9R�q���;���[��n<�sʅ���Ѵ$Fy�cxONL��%��tm�kpa��y��Ͼ�b�#(9ϯ���]�����hm4<�|&�s��=\��2~	/�Y�-�zaP�j�K��������/X����i���k[J�����2{����c#��;�ze:?~qи:Tц���H�W~�U���&���jɜ%�{��Մʠr��o���{~H��u/�������Ջs74&<Sx�T��Tl&�/P���ԼyT y�D�d/$��(Md�P��9�|c=��(�@��"�����8m��-?bp�R�ƞfּ�~�|!}[�aub4�WH4w	!Φ��è�QaK�,�h����y��)�1H�]2�-=Ad8<��f����m���`Z
�T tt�����J����^���~,�pHP��źb�`�n�ry�pE�����!�}\T�B[�#z�y	��Ո���εW	�N)4$��@�����<�64�X�0��4Z[�F�7ɯ�/��[��wRoT�g��~��%����1@���L����?�\EPd�f����K��C#��:M��f�u�`�>��=D&7D��^���;Ң}�+t(_�o�I"��2K@ST S��h|1��e�9��.w�3	 I�e*�Ю2���1S�L�F�t҈8kݎ�9���}�O�W���ZzR��pW���.���X��T·9��-��&E�Mܣ����/�x�2��?�S[������j}0'����Z���B�*(+&���J%p(��20�Y��m��k�5��� z-�K�T@��p{^v�9Wx5vA'3�� >*d�o&�8��Y�wU���.�B���j\����R&.�9r=�l�=_1A�fJwD��y(Er|j�H����٭�����p!��zב�kĹYuu�����6�;U��.�;I�w�D���7t+6sl[ �t�Af຋�N�����Q�Ȥ�E{���w_����{b�-U�g�џ�9�R�w���-�L纉|��_s��;2��O����<<`���TԚsz�A�*�qu�D�B�?�*h���`k]���ײ �k~u+K#n>����>�AJDM�ί�>�<�,��OP�e69�� �7"�ݙ��奚�Y���swy�- ���#�	�e�zQ̬�����f�g��-9^	��dt�nD����!x �89���W�¹iz834y�@Z�'�!��m����r����C\4�	�6��[�U]�c�+쾽�a�+.��_�7u��Eʅ�!��{�e1]_�]�G�uv,F�3��R�C�8�?�f`�⴨W�Ck�\�����pX�!�la/v�2����G�ћ�gy�v�K�����w;�ZN��2j ��J��k�%;5�t����I"�W��h�k-P��2�5�u�M�\����k�����ɷs�])@�����Š��>�7� �ɛrǊi��Q����*�0�`<)��B���(<�i7�
��Rw��o-<'��v�Y���xӲ%�*')$�f�b�s��nEi��Vi��?M�r��Om��� /�yG�%$�p_ ��2l���D�Xg��B�՝[�i�@y�Tp�Y���(��]F/�ǒu�%U3)�σB�ן�^���\��ب��jQ��쓪
�
��V<�wɌYϤNsf]>�#o�O��e�dm�O����e�,���u(��L|��=��㮨�Þ�
�����lEr [1�%��1��M�e�o�2v8ɺ�*e7pQۋF�m�@���.f�'�eF	yƜ�7�;Y���Y<�0�������C��y��s���c�UȨq̧���� &]G�k(9єs7��(�F�N�6���d1����s6o�Ch"`U�,�����!�ymM@��\�'��I�{*�3���?����	�����&HYX��z�A/>�|X�Y	2�HEN��a[.�c�Y-J �w�7�n�C&�<��?O��-9���4
9���a� �U��P���L��t~س� =��{}^��ض �ie:�o.��N��{_2���ۮ�uPҽ}j�׬$���/��������֠݊N���J���j5ZY�v�G��.��J�,���ed���j��� 	>}���"	��}|BΖ������n�QLy�t �%�AH5���.qZ*�S�����-p����g�����g)?W���j��M\�)��Z$xf�C��[��N�Y��	���n�y�����+,)��'�Ӱ`=g8D�E)AI�F�Fl��i�ᵸO<��0p�I�V��Y��e��d���߬��9�FɆ��ьw�[ROoR�����������Pp�6�׿l�ԙ���-��Ű�r"�	Ƽ}�@�&*��uɂh���g�99F �����f� ��Hc	剽�3ߪ��o��kf6X|gi\O�tܰM��9���t�K_��Oc��q�vC���[F��k�r��6�:j��	7�*�K?��Iv���m�bX�!��!�"��	�n��3�<��F'�(��(XC�+��c����lu�E�c�2F+J�
z�l�Y��ө�D��[��w���.79\�o����EZ��p������������@�����#�RmM�P���᪛����V�8)��֬�S �&�c�X&�f2[AB��gN�(�yˏ�L.��!�ALa�w~3���)����36 yȠ�U�5��зt�6�pS��tn�s�%rx�DJ��w��ꄸ���iy�(9�{ܽ�
7��R�`�S���-�W�.����\�Տ����Q��"���ô�*���Fk��Z\(\7j	�0!4?�`8�H>Ң���۵g�Ϧϴ3� �Ӗ:I+L��tjk��T�1���4��H�I�O	�8B�-���qu��uPo�����Z�jL��=���S��%y���hվ3N�o,�i���.-��ip@���U:&�>�>�G�
�V_�ca����߹�W^R���߰ŗ���ܰi%.��bS��ޜ��C�Z��Ii��LbLv<�l�ۤInx �[�^�L/�~4�^9�{�$�#^X�aZ}%�_�L
�USr��~Z�Hv6���)�y����5��x�L6�|��}G�֔nw?�s�"��<V����8Nn����Hl)��Iͮ�\T.�?��x��ꮸ�6��A���}��a�(�0g�J�jG|�� �I�4�������_� Ѡʎ^EV�4�)�Q�I��V�%	$\ޤ�&�}_�^��n���k2���i��ʰ2��gB��j�~ S<m�
���x�_}I6��x^��K�p��h�E(3����&��fY�12} %�9��At��T�1��#��fok�x��z�JG�V^��83Bn�+��o��IF����~G
�$Y�����Р�*��z��⟲;Zip�}�BPp�W�Q1�E�r��q�a0�%Z�1�%t]ړ���u۩}||P��kZ���1��7,ޠjYІZ3���U��Z?$b�[C�v����7�!P;�?ǿ"n��}alϾ������wI�˜m�{��E`�B�M��X�Z%쁣���ڨU��I�Ŏ��CCC5 �/�4���c`?�h{�a�A|�B�'��}�
}Z�S�+e�&���{��3�|�:����2I������7ȓ��m0��a��
��-z�mZB�[(��qIO2��e���8� ����O'qQk��m��"�n�(bAv5Ct�v�:��n�1K����NP���"�TAj���`�.рr���؟P��j�R?2�a껕AsYb�����h�L�s(���_�8�<?o>�C�BJ��w�M{=>@k�;��m�о��K����%����1�'J����J=�Uu���ϋ��Ǌ�����]��${��J�q/D|-�P<H1`�	ɓ|�uG��Dr� o;K���£�+��0��ܿo~��)z)"%{=���%W�mԥ��-������8�'"n�?��a��)��d���c�4�[Х�Q:�?�JRw� ����rK��~�L��ݹ\��GT��c�"JTO+DlJ��?*]�t�C_dM.���#��$~a#ȸ{?�	{u=0��[�៴� ~O�2��j�.��3�z��=�2/��_�ػ�c���Y������j�᠂�ɸ���W7Y�U�,�cX�� ��_�,�x�ř���[��U$�gԤ����V�Dn#̜K���w�0Jy�����C��v�zûE�h�1u�#���T����F��$�P�!;���,�zLΩw��x�J?���9�i���0�i�.��)��cUk���,ЧYN0����]��ۢ;Z!�Q�L"�R�#W��G�o��)��+�Q� �G�\g�)f6I�T�6A'��	�n�L�`K��DL GFZI�M^w�z��uZQ �I���!Mp$�U��C�vgt���vh,�a��7�¸��WV��}��R8��.������i�C|���>�h3Z�U��5k#���q�4������&���J�y�ÀO�<�^���� uE�6tH�� 0�{��$&b�@�>�2���V.�����m[�.����+�S��|�V���P���սV�,j�c Tnb��U�0(=���si g��9ܰ����9J��sȫ�S��I��ãn�/�-�����A�L������Z���Z�'J�O��"GZ�q~&ꙡ���0e<��};�](�T����u.�z����6�P�8��@��1ao�&Z�P)�*ϗW}�J-���w��?Ë�;[$Y�M#I`�ĭ!�m�ħ:���J���I�66W`S��+�27�^����"ڧ��������F�W�/)|��4��SZ�]W��gx($�9{,7�����3���U`��"��0b/��U9�I��k�/��A���6Y0�[;+���Fm�rHtYwѠ z��2�h���(c�gٹ�v�Վ�D�
�$�O�M�N��c�gcy�������m��k�!$�GDJ��0cؓq�e�: lTo޼��*���-�cA<�J:����	�AKn�/W�D&O�y����$J���L���/��+UMٯ�z-$��)^G)�PW���jl��2揸]��v�@�o>>�5���I��!��u�V-6U{#�[o㠌��;�-��`���1m���Ag���5W(�#PF�Z��`��3uR�E�rI<��r�$XlP���t4���V�Dw��	v�l��>g���r(�ٟ&�Z�8����Eq��=���P<��=[�h��LR��o�D�qV�3�ތR�[�j\s9�- -ԭ#e��J���M���gF�s����q�C��r��K��oáHv�D��&�7yʀ^5#&���Z�폥�~���C�;V�%��
FQ�<0�u���2��)����ټ���K��T��P\�xH�	4��L�7��R�c]I��t	�؋_<��Ĭ�ޤ�̸2\�?h=��� !f��ӿ�Nx�g��ݿ��*BИ|�ed��r��6T��Ԓ��;����S".�f܌�n�iB�^^��`:�]z`l���F�! 2��(�Hy�'Y�=v{gÏ��k2j��[�5n�����Q=�ŗ��Ae-$��dT�� 'x�u���)p����"�������|�Vǌa�'߭���"���>�Ѧ1�) [_���ɣk$Į�x0��}�lH��(t�4���W7���~OZl��ԭ�D�����[(
gg����i�4���(��vm���k�vӗ�)'���pɕ�Bٶ�;��}+��AK��[(D9>�Wy�֕vy���ba����,6�}�7#[`���Ak�_��_����1G�j���Wȳ�*M��\~c�I�@��N�J��5r�2�(\�	�8�8���nMxX)�(�4�H�.*K��CT�0B� J;���$���0ԍ����G
}�rA�V�����Y�]���2y�:0[!~�ʕ������ �E1�9�E��2�0����=�'z_U̗��)���=/���m@F��r�/����X27f�	p1�A�#>q�YN�?뽻:����Aţ�W>Y#ci]�l@=2�}̚��m��~$�����=%��,F������iU���<���uW��A�}b����l�D�2����}�It�x�q!��U���ZV}��Z���y�wT�Q"���p[�V���p
�k24N��aok*s��Mi�sW��t��`r�re�p�Ɠ���@�< N��.�^��q,iZFWqD�h(��1��Oӂf҂��tX�Ѵ�Y�6l�W�oԡ�YV�6J���t��Rh��������M-%H*W+����Mb�Q�&��	��D#\l�=i�7��������sj	�\��U�d���=���.�
WD�z�SY|Z�\u���Cp�ġ�����!Ry,(��vF4Y�V��^�8�S��"�{P���(���̍�R	��s�`�_oC�N@�I������M��t\�}3ű�C�"��p����1��a84�N���^P��@��.B�4�g�3c0����1��*�TƦj����j$�v�}���W���Q��hNU��-�>;;��H�{_Ω(��diGq¤��jWM-�>8��'���ֿY���6Y���/ʺ{d�Ȅ����2�pD��L5U�"/ܗ�X��xN	^b����k@�g�:��%��a����XC���q&%	�����ME�閞�8�)]�5�����Y��{��{���	�p�*��a���6))u��F\��t@(�op�D`y����-���v
�-�����l�y吴w}<s�z�|�%���P�7�^�G��Ԋ�t�y�C���ƚ�E\�#��Q^�;C��m��:�(L�{<#���#*�x]���k�e˫�E�J�7�Z>���'q�H��l4�-C�]����a?�*K1:i�^�EvLx<y��v��v���TM>@Cn]�M�
�纱�O �W��`���)'�K��kN�J��]j\r1Ehշ~��$�-�ޅXU8U$�b��q5w�輳͏��_������r(_�.�Jr�Yǘ���?����c,3��]���8إ�9�M�Ut J���YY��!L�Ձ�L�]��u��I�ӐJ���(�إ ���g�&���zCb���]j5֐:�KD�F^Vu�&�������Q5᪪�yod���%���W�Ne������4��2,��fw��Sdi���w��$�������+�Df@�ކ�}�gR���@oS��3�)/u�`�,'��%Tg��+��~c�E��b	rs\�����˒�#L%*�BLA֯���؍�(���"N��e1����TGN���8l�P�����j�fEz?��H\�I�s�o�fq<�W`E\�Iɝ<��U���l�5�V~�22���hmac�1�.N��mhѰ.aj�$��)܍=ų�'銽�"l�����l���3&/�����n=�r�S_i�[_@s �Ǖd�nFL���/��j�Y��g���Py���������S�4J�9�n���|X�FR{,�ͨz�����ꖳ�z� ��Y~� }�SkY���L��%2X-�,f�=���j[��6����_Vh�c&�m���+	g�]�N���y0p��$W�Q։�����9��F�ȝ���Q����?5�Hp�ϻE6!w=I�v	ê��v{
����/X�4yc2b�?6ԫm����]�2m��&rM~���X��zVh&1�Tc�J�xx�y[+�L+7��5r�W[���M�]�D����𶋱�����lEU	ЂZ��õ]����x6h���g��8��ċp3Q��{��fH؞4��+�D��_���;C���d�l���X��:�{H{YM^�f�*��� ��V>g6ˆ���8>s}��sZ\��)�v~�kd�Z���<�iMA���n4�7�����4�杰� E��ٴp��3��G�S�� ���v���ng�R}a��hGsg&*�6o�����i���UL2|?1�~�D���%�k�U�zVKŧ��:!�ڎ�L��V)ͮ��LfI���-�rG���i4�>Paɒn�J	[A���Sܑ�>�#�>⧟jG���b�5r�$l�Y�X�⮈z��
�ߴH�\��{���y�o�Z8e9���/�b3ea�&��B��l�ea��_�+�!�."N�(\ �.?l>���b���4���u��7=ıu�0�x4�C�=!^:��B7���EC�]zD;�To��#�$l�uT����i/�(#��Xܦ���l^l����䢰�����^[_��Z21�$.��O�[�IH_�{�N�h8��u�Pe>����Ʊ�s�=+^����35gn���Z��{^d�~w`ȄKWH&�l��<����x���{���k~Y��d(�:��v�w��rרM	���0��zQ5:2��eч�C��=���Σ_�l�|O�Lu�#w߅��c&=�o��k�"9��/ku���=⚧��(ƌ��~*[�����* ����U�y�	�q�0ɮ��^�z.�m��蒉8̽���@*i��W�ns�U��%83�lbl�'��3�K?7��|ւ	������f����W_#X�~8��P�dI[kGqūh��5�6���R�H/X�9�G6;�֐�t4�١!�p�^p�u�<�= j!Q�c�����5���(e8�����咩`�����N�[���A�*cY_!��ᶅ@m-=��ym'�}8i38`d4ѱ���F�kC�MI��xS��}ziw�콎	:<�-L�[X�想��V�)~s#W俁?ozn������e�"�z�+ �9��Sau�.��
"7G�N �C���/�`h�QP�+��h<3�I���j��
����=��������EhƎ9�2��H)a��σ�����z�ΑN�*� �%A��0��,�wWX��# tCG7e4N�\q�Q1va��f�j��~��s�J'kʤ�Z�Eʮb(�^TL�0,��gO��൅��Ww�׏C�r��ZB:�l5��hbG����)��Hp֍��v�E#H*c%�V~n�D#��l[)�m�
��6K�=�Ě*��==w~L��y!�R����^��-ύ"� ��F��UPJWBQ�����0t~�'�mR��C�vP���'��"Q	;8����a:�7GEa��
�#H&2��q�{*h:�!/_��ȜgF�HY�F�nn�m+��}��5��,�#S��p������}^�1e��>�gʧf��xb"��0�l�ĕl�}W�Ŋ�U]����u S�C��f�O�ѫGgR���=b��*�v��gF�KׇeE�����p����B���_f�
��f�e��-b+�̦�kSom����
�=�Z$f�x�����z��zn�3�P����?�mE�f4ڱg�|�/���&[h!e"`��2��u��"���VSL2_ys�۸["Ϧ��.R|V�*�����@dw=u�Z�n��6�?�[a+6'`cF�������HK�p���q0N�)v�7���@�G(���2�@�{Vj�=�T�hO��U�D��9�Hˀr{s#��/���0Rk��R�����@���4-~���ʷ���N�֛��n�piK����|^oe�Uv�y�H�ʘ��G��p��y�q������\�k.@uo�qs�c�y����54���K0j�h�@B������}P�ԍ�̟�h��JݩTsgIو~b�2e{% ��n��-_W~J��b/�V@1On��<\�51���0�Io/:(�vM�]��s������3֠�?�t��0��ۄO$S2�[�JWj���}D��3���Վ;�6�p��N���	N����I����(Šケ�p7ۖ����mq�Bq������u�0�3�����EY�>�⦯��+\�th��d�Dܪs��p�:����<�J0VFq���D���veZ���*ID�1	�n��h�ռ�mĄn�XHH���PꍝM<��"�%��4�H��d&��x��;T���O��g�j���>CM�ē�١t]���9
>�Tg����5E�?&_�8����8�2���W�R�ϻ6��Z�"�k�"����ob�4��I$�Yi�=B&N ��%Rv�)�W�Q�T�}er�F]�g�S��z�-"����둮P���":�I� S�Hb:����ޕ��I��~���L�u�����o�Xh宂��^����\!=ǂ���$M��e����5�X�>�飏w�tg�����t���W��D�Hh��D����S��O�p���ae�g_�C��F���:�@	���s"R�~W����ˡ����'Y0����^��@�9=��G��[�T�Ŝ� j&\�ׁ�	�	�f��L^GWg�O����h--�'���޷<4*�#:6��b�YU���`3���䣁];D0W��a��ʠ<p�!����&��Oi��W�"O��V�ʾ<����;��)/���8Z=�%il4~q�n��X��>���J|�3�$+�Է_��F�J^k#��x�/
� A>�$N)dܿ�>w� ��8Y���|�jߡӮn�|2�3��w������,n���:�k�o�Fvb�ɁDHE�)u�M���`��d��h�آ;#�J�[�N�a �fI�U g�����Gʮ��z�!����_��2o0�Zї؟����`Rɶ�A��	(x�"�J9V��1��=(7����o���<���4t����t^�%h�ϐ{?�9�U��閕;ao"����Iݙ����[M-�gzx��T���2�%�� �r
�4�K�S9��]^5�3j �n��I�%����o��d71��پ(�֎��}L�ٰ�/[Me�%7c��9�L��!B��7 0?�[�c���X`��ث>$����47�+G�:z���le��a���<�2���uxpI���&�9Ң�T��}3����PB�IW�b���TH��Bgt�l��c;�f]In]<;ш$BAy<�O�ύΏ��2�H$Z�W"�Q�[ʄ�PPs���}�R}��H�Tڀ猋zj�y����|3}ʈ.~ =>�X}���>'!]���Qn��m��SS�����;S���S�+��i��wax`�X}Q�V� ��o��z��8	�f�Z{���-7�޾�̟���������ⲍ�,&a�v�׵2�6�69{��r���}ۅ�<KA�7>vn��ȳ\��������
�#0Y�<7d"ԑ�S��f:�h�L��E4}��uʐ ���i���b{"(���'�R���j�O�{���`��H3��X;�#Pۮl�=���]|��,���ܢ�-$���;�9U�U]�Lk����d���-�����_b��}���ʄ��KC�����k�,��xunN�H*��o=��[)|�S�V8N3TFs���挛p�:Bv,'n���r����@���DMk��NG����3d1�W3��=���G!������ )ӌ8k"[���m�ݳS�ģ����������ij=-3䒟��Zv�Nq 	�L��������;��Fl�sqj(��^��:X���a��|�VBA�!�\c����E�OF���X n��߼-�����r��.5�ᘆ�w�����^{�ӛ���/pǄQ��}D�T1 
ۡ�g��T%w%�?��/�P��6���3z���Ғ��t��|��O�%��@a��*��A��P�;���B�­�B.�_wr�<:���Iz��ߖ{H�R5����H����u�nn��p�I��=V��Tq�鲅�V,uIan�vD0�"���
U M̨����JJ{bJ���,g�Z)����GBP#{PE��#9J�xY��@�����~�fM+��}��z�����K�Âfޡ?�!?b�d�[@D,��n�@�J�7�ʖ;g��9�
��ҢMb��f>^�����?К}H��x��iK���w�����d�=��*ׅ���G�W!A���t�� �E�cL��ڳ��J��@��U��hg���*� H���}�����K�D�6}�.i��o07�3��i�i�Rޮ7��^..@��?~3pb �0
�gA�:x������`b*u��&鷏��8�q��
t��o���\�����d.�t�]�+� `'��2�i"�y�����p����yd*�I[5H����@�S�Q ����;2�|�v�0��i��=Q$$_އ#��B��Ýa��Kp�[B�0��g��L0��㰣Ï&�e����H��N�z���q&�2A�pB�e(?	�hۑ�c��6�i�t ���A�[�v����?N�;����qz_RS��8	��~�-�>	�9x�WGf�ң>Wja��p0�OױZ 6��VP�ۧ�c	B'�>�ߊ���
��k�)����Gι���"'�����8���w�9˼ۚzQŬ;�pE��c�m8y�f��^_I�K*h�S�+_��3^�^�����F�G_��s�'�3�z�E���{閂:lhD���
�vTw�Z%9�(�8l[�i
I�pSH*�o���&���B!r?lZ�X��ԩoZ�����Q����&)$�E��������!Dy7={�w��Ύ#�A�2��U�l̚�t�L�CO_u7�	�ޞ�Ɂ\�%�PU�<N��,'���^��ǣ�&�>��I�n6�}R7[7x��S�,DD׆�����D�����&|����$I$�	A���|��Ap�R��tgQ�>���<��k��63�=Bce�ۺ9�����?Ӟ;�`����A�))
��?g.L/�2��i����C��+Ә�i=�Q����*},��??E��AeRs/!��@��4���RU��gSX�}����R�]��A��E�b��2�&�ܬ�!�^Y$����1���g
�� �k;D~��9��٤�ښ7l�V|JMi[^�|�w��ks�>��hY(�-H���Ѣ��pz��B�X'�]n���WB2/�n��B���K��B �#��I%�<�R���&�h�+���C��4�����W[��'�O
�T��5����@e��m�~%=P� �Y�vuNN1�T�s����(��lH�V��Ń�L#�V�C1b-��}bx����? ��I���ؼ�E̶itB�|��(ǖ*~:ZU��,c�|��=:�^Z g?�+HzP�kʨTY Ah�&@9M����0���C�:�4��>a�e�,٠ۼ�ll�+^��5�B0����F7�5�KX�ۈ�b�L�I��FК�"��&�Pچ.�����U��B	�#Q�FD��Yb���˞9���Gl����^yUX��>��U�!�$�c�\���K.FZ��M:S��OV�H̃�)��ڗ�<~����
M���S�\�mOMx��ύ����V1z�w����� N�'֍U%"�ڄaޱ�!	K}�  �D²��s�feZ������~W�T�K�r�C] 9��]Ex}mC�Bs�v�қ�jm�n�feM����N7���T��7tqϧ<9g��vH(`c�`��ݎP]׼zpH�����%2�$N�X�\q[j�O�JDd�3���%��������r���.N����u�4��oxV���|�|k�u�Pe%�$4��o�<0����8�5����
K�����G� ��yUa���]
�|��p���?T�3A� �Z3-��3�#'�CO��=��������
��2�]'�SFE�7�_b}�ܮ�"�.�s�/3��s�cv�|����?^��vM�.������WB���ڣC_k��O�tL��L��y�ĸZ(/�~�j� ��2p�b����g����T`8ߗD��U�gMa�$n~1�D�45��.��Y�@�&0Y�#6炃T��q���L���;��k5K�B���ܘ?�!w��E�{�.� 5q��7��:X���1<x�Q�^���J\$z����:P��:LU��kg�Ĵ��n�^�Q���6��2ieJ~��^C�D
+3[G.�	,�{��,_T���"Xգ/�(�!-)��*��܇��Zܢ�Z��ה���u���j�G���(����.�k��G/a�瑟,�I�Q�q���"n�g8�����H)��4�(B��s}ַ��,=��Z�B��FY^�h�{�Sh�\eR���0��MaV��>ކ 2�5�L�i�F��@��l��(�F��u��A�nn8�Cl�N{'q�P�e��%t�j���C�17���zDq�Mu�'��Mٽ��&���qm�v�w5#�}�H�������q������ފ�t��2į���p��/���,ȶ�����f�9y�B(�0�C��Nn|B�aN3�]=��)ߙN����>��jIz}u�J��]F�w�����=Dr�{�ގ��눁P��1Nl���������k�Q>;�3�G}�2MI��4�$���z���#��08o��4�g�Mh�.e���Xr�*\�f���8aA`fa٘�\��(�t�qF�6��
��06�S�:���Z4<��ٷ�X4���l��C�~fA�:�&3muB�(_8�W���H�Z܅�	G	�e��U��!g��w����[����ikl� %��C�P臺	�9���=9��ٯ�/�!�w�t�&���򧈦��`9��8:��D�R/�����~�����		O�`�+���{�1m ��ޔ�F~?Z��1���	T3���%6����L����d6l�0F�t$��:$;�rv(x\8����������:��С�!]�i��	�>f�~�Y%�y�hN6����u���p9�ݾ�\����_H�	p���m5�c�d"iO� �-$�Ԟ`�ZAF,l�ΐ�h^z<���b�zv5R=�Z�q���i�~�v>���3�H��L)�\4�з ��^�b��bcj�����t�h]������"�z�T��/��=u{��S�[��F����M��p��}�k�EU��.T��hY=�H4*G7T��ƐM�Uh �XT��<nV�^��o?�=g���6z��gu�ou����5J�< oV���Ki[�e�Ѡ���1W���
[Ǚүj��aN�h����n��.B�P�����,�ɭI"2�u��F!����	G�|�[��ݗ,�WعXx�}�����`��*���X��MB�;P��Uȫe�E����F�#�e\'$MA�Jn�r�8z=�7�k���O���@��V�L�Q�$FJ���hT�v�3I��1�|f������8>��	%�t�֥;n�7��EӒ�t�\u�U���n2X�g�=V�=œVj ���d����X
ߔ�>�6LӉ��W|���$j�^:�\ o/�ݞȾi��>i'ڊdG����pW~����e�Ij��l@��.)�� BP-��oJ[}�9	�� �
ɺڕ�`ŹfI,�P����`&plTS�zW��ad�|F�lsl;Y�~�A35)b�B�5Խ�V"Y}t���ܚ�����5�B��F�ޡ��EԮ�c�x�i���������%�T�RT7 :LCK����5ä��r���`/	�Qh��S^����Pk/��z��㲕<��[�,����sd�����;<vn���5:%��Y�J{�pf����XY8����BHueA�X=�s�Ķ�I~bI��竸2�J��/l�T������;`L;����\(
2&��T6�@��
�
U�"US"�w���[������\eksac耴�}�cGl]�͘���:/���r^�A6���{h�tj�p��xw�U)��F��C<3�'�p��v-�e'��oK�O�J���c�d:?6]Kl��wO8ǋɟ���;ܑ,k�h��5�77�t8C��K�-V�|ē�˅�㱱M�%M[� �ݢ�&(K���QM�֔���Q@;{^�!�����*&�f���g�s�+��\9��*z	��g,���%��{8�kvS���+⇻��Q��B����jn�@�,���R�m|^!�}�෉'���grp��N5L~R{�hZ��]�_+���!��.���F�`�9��12�NW�������q��6w}��@[�T���Oo�esq��ߧ�KMe�sUС����"��Br�zq8��{������wańi�)�l��x�� �r�����	�������;
pY+e#�R�~I�h|6�&�j�$6�9�-����x�Q�^�V��e�"�"m8��k K��dM�`W*3n��2
m��J��hX���������+X��7��*W�Yݺ����F�
\��hR����ͮ��Ls\��v��P��bK<��q�N!/昼�*���8oQv·���u�"|�=\*�#�ǰ@����&��)�H�m7�0G�>�Wb���{��H7�$���0/�X>a��b����]���x�SO�z@��U�٢ŏ��q�o���"��tH[Ѩ�=]B������-�Ӳ4�4xY�"sp��Β�5D�����G��J�*�"?M�t�pt*&J9M��d!���[�N�2��i��A�8H��,7%�>�A�ce "�䬸6�9�Bz�z�ccB�C	���Ų��� _��3���(�臂�<�]���>�����̄y�cL���D��>���;����J���9ovG����l�<�G���7I� \�۾�#gu&ĸ�&wg�m�vp�*���=�X�ҷw�ܽ."�����9M���c3Y+�p��sh8!F��� ����>uyk�*jE��T�ف6ؠ��S��{��?��0{,�wd���p��^z�����j����O�����C[�����O[Nu��M�M��'"�q�	�gm�#ښ�f�ͦ~m��	&ݸ��Y��{ӓ<U��A��|�j>�͔)î�<w^��UT'S��Hh��l�7o�����J�ֺ{��K�Y� �$�)d����:h6n*�m����8�l�]��JV&ٓ�g����]^ֈ��gG��q��bB���TWzC����f8��O����5-ة,4���T.-4�C��1UPc�*�3���o�P>�B���r�ۂ�)�Y*9��7�6K�Y���ޜX���u�;�¶�R���&����B���9���v�f4�_e����P��;x�}�,�x"�U٦'�\�-��y���ko�ۋ@���9�Ay'�:�2ŃB7Gq���bX����ֺ|�@[��g�魓x�sZ;��#�5�H�����&ʡd��l؞�����;Q�i,��U�RR�t��[n7��b�D͜DNk��J�< ]�Կ��䑾a+t������b ���,�NT�M/��T��A�c�}�=����)�(����O���Ff��VU��6iI�L�c�b�>�%��U>�����T�q�h?�pm"��v*Pc��u}�5N�j�����Q$����i�:��䤲N��ő[�lЇ�����R�$o�*čP\���#��Oe#����+م�޸�˃����`-gwf�<�`�� �	�