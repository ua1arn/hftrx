��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b��K�G���Wp����&�7�����F/7�,�9R7.�h�r8�G{��~'}�<���7�y�<j$��6q�=O�NXb� �-؇X %�,�ԯ��� ����S�h�떋�Y�M���� MYo���s�����.�a+fy��r��0W��Wwx-�s
��b�A���b����`��K��/��ٛ�B�o]�����=���a=+ �g�뢢��a�a�$�ǁr[�3��5D��k?��a![�K�F@�'x��_�o���~c���'mf�]θ(�K��%�c����^�'��»�jZ�Oɉ�q�'L߀�	��al�>�"�p�n�}�7�a9�4dH��bEy�$=��Il��
3�X�{
F�c���. I�h�&��'h���w��|F6gDc ��	J.��֠S`�����J�4rl��`�s��td�/���F-��_ o����;1�pP34��s]B|������au�@�[^��;�ưb�;<�Y��LP͂/D]�V��n��W5�Y�̴	���� ��k��{�,�j���.����Y��!�4�=1�X�YghLOof���M��L�}󦰦��0D��볕6����o*�%6������C~~�tP酁��mr��k.��. ���Ǹ"�Cf��aIH��d���jO���ɤ�G����-R@���}�mV�2�vbv��o��e�ʒ��_����22#%Λ"��jR���ܯuHta��i����V�"�2j���g���O�ª�p�M�����������Z��70�����BznA�/롪�l#�ǧ�����5\4FYOﭞ]6be�����A޸~ޓC-��ʚ�k�9�P�˶����J�&Ǥ6�R�$ދr�F��ڳ�w;��S�UK]�>
ᮼ'�i��%�L�k�$)�3������U�O�.�l+8{ID)�����+��<��1W�h�ܝϛ��N�݈3���pnG��;&HF��5}<[T~.��{*f��da�j�}Hz��K��"L��y\��Wб����"�ox��>���+~�.;
��%��>�+Ϳ���-n����)RXR���=����3.ʧ)Y�<3�w�͠���r�]YQ1Ac0@�NX���U��`l2K����f���c`2�A���h��1X��d����3)c��|G��ӛ|�%"ds���[A���
{i/|�ɭ1oN|#\�KR���P��y�6���c�@�V�s<��\�x����+�Z�]���ԋ���B5lм'�G��_�?�l�S��������q�C�����PV ::#�$��6s�@�;-��%۳�]����b���'.9fR&�B���_" t��<1��|���sR�ҝA���,n���B��%i�y<�$�a���!�6�ۤf����11���_99�}�LC�zivj� ZMt�W�2�m�p/����}E=��.�)�j�C�i�n[��JgC�͏`��P�ڙE��e�d������6gSb����<3��!�1�1"R]��]h\}�-Zd������|�t@�=mc�Z���x���8���'�o���Gx��ƈ���6K/�}��Us�+�e�V���Q�������3}��K0<��稹�4�����������fģt����c�]�I�)��'(/�+/u�]�I�(9��@��8�(�R0m���v���S��2���ˬA/#$^{��[�f
qM�wz�ů���O���vi�������NaC�쟃�N>#�c~W��c�	��@�s�f���s,�*b�{�rlt\ši\Up�1yE�	����l�h8��jL�6[�Md��c��/)^����cjNH���&�D�d(��#E끸ڈ�Bw�2 �EM�l�O����R�5v�A�f��� .��c�"�_�}ċi�:���ʎaꡪ�R�<��z�
�g����٩����n��������i��JZV�I�������GR������#c4Bs'+"����ˈ�8݆C����ӽ � �=��1�V4R�8B�,�Z��]A�P>"-.yv�U�}�z��.�M��<�v�!1gw!a�fQ�
�.롘>�x�X�b�g, _Hq:��V��r��e���-�<>M�H[�w-�=�H����3rrlW|Ju�<0��������ŀ�Je�Q��imW0�_�ʸ��$�-Z.+�\���!�_W��@h\����]�2W�0�|L_��vOXJ�&�o�L����.f���LM��!�V�;a��gp�
���v��^<�`{�����Ky�|���ɓ��'SUyih�[��:(5y2��"��Ln9�m⑏2"��bCb>��a��z��i�k��(E&����U�<6�Z)~:W��:̡^ǧN�.'0U�xJ�r7S�;�Dώ�6w�}��hc;�����}��В=ֈV�h��:2l2�0Ïg*u�饙A��kUZc�{֦z���	��#���FE��=h�o՘}�(l�#>?��*�bE�V�yl9�n�x7���[R/����p�2���̐�8����vF�ZQ�0}e��.!�����a���*�\�/�Lv�E�^M�b\�w�S�����J�K�xE�E]�n_%g���-溫������HR��B�v�@ S#��+A1�Z���ơf
�V��K�{������~~�ht�>��f�L�X\ٲ8�{��&N���:��K���w���0{���q�!o\{�Y��U'�ݖm����,�1 fAhө�f�� zL-f"F���.�����w������� ���2�N�?�i��W��E���_�	%"l[aH�J�1	�5t^��0Xߎ�i0�۶*�M�D�T�2o	������l�_���p'#�&C�ߛ�:T[gyV�D�2o�6*eК8Ӻz�X���5��B��@a?qua��C�^����n\��_Z��^��E�m	@��2E��F֛�k`�<*��ܤꍕ' ��=���#$�R�]@����7�b�q͟VY�(���^獐=�y(GƓ3U\u���'�����0�nb�6���`��TT|XX��yҏd��Hx-��)�1����|S��4G٤94�eE�ڎ�'X�Zm�]$/��9ng��n��.[gH�S�K�+���l��UJ6+�AV[do�ֈ@[-,������GjT��1q+4��t�`�TP��z��K{T=m��KO�D��ϯ��:�
�� �x%�rs��3��	]_����.��03�eqH�J/���(. �[ˋ�%$�s|�z��K�p�K�����ɸw�����Å�PQ�b�����G7�֓���}A"�4g�=�'u�i2O !��:K��H�ю���)әQ�߇�6˦���v6$��D|!b�}�A2߸1g��"�w����Q����N]����JjEߤb�E��j���eO=V��,���>`58`������p���C���!���N�C|_��:
柈� G��'[�\��a˖%�e5����^�@��~�<Z����O���~b8PR�Y}���������|�y0�5A��囎s�g�'���JA��N��@���緵���-�;���j2�هI�<��yѷ�%Y�~����T@h�~;�R-;#Q��.�����d�����y�����P#o�M��\��Q¯��F�Z2զiA�w2���wp[�����Ͻ$;�Dv���~��x�Bta������=5�ݣVz�I����C�\ܫF�gÁ���ș�l�G\�Tw@�&�d���U�,6�@]GFۨ��0���YMA_(aw���3Mb�L��c����v�L����ħ�e�4L3m��q�$��V5���G2<C�N�IaG@eM��S��A{TL�r��w}χ0C ݡ������כf�H�GV{�ݐ"�n^@2޵9u��/��J�uۏ�=De5�DЛ�IpH�iFİ��o.5RO):m�3�F��Bx����x�&�"���e^h�r,�8����_���{�_"����|��4�`D�d��w���N���j%~]�1���ʾ�&�dv��-�ܻ�$(�'���ݦ�\�g��i=�e�.�H3n=E�1t�s&��jЭ-���%�fO�u��e�"o�X�y^Z��P��M0Q��om�����hWc��l��!����}��ޱ��	�K�����'�v���8��M��^)��ҫ4�>���]˘Ä��zq@X��tLXw��]ɑ+y������\��1�((G^�C/5n��Gs��nwb���i����<�9�~Α"L1����e�C�i ����X1��DKa+�Ɵ���{o\���{��Q�܃�ՠ�'�%�A���+5�M�⃵6� ק�����p��[����a�������*�~(��$)�w�;Q��	}����^U�$��z�8�	��Ŝ�Z�4�jj�k�G=��̤����$n����iV��][�ܫ70����HM�k ��Ąatm����C#�8�B���?te��}�v%�̃d�\����k�+
� �Z{�������SfK�<�jI�@�6F�����x�Pw�|͵��-����,ǛA�3f��}�t�7~Rĺ�i`��ȯ�Mw~M�y�p4�m*��?+7� �8*���p{��ɑ�ǈ��GU˓�j��nm7qwW;(Us���+�R��g���iE��P�Q�|[��R��2J�|�L8�-1�ȍ(�_=�Ȉ�x��̂�6��}3x[�����浹��DBB`���R��t�q�s.�^��B�4o�ʦh"�$��U�2���޸H�(���++0ć��� ���?���C���9�.6��yC����U�S��#�6e��w�G�|>���˶�Q	+���nuS,9,2��Ϛ�7R7s�Hϩ���fau4�d�F�g����{"9Pd�&�^2|Gv�ic�ul�Zݚ����7�⬈��G`sD}_������{j2��ڦZ�ׄZ����!�J�Q���c>�p��V&���ݞ��m^�T(7ص�d�mk��V���}��b��Eq���Q:p�l�M%6Њ��a�T�1Չ�T?�EB��K��$�:��uEp�	��q���?iOT��-�(C���� s G7	�&H����� �[�[�,Ɖ*�Vʂ��u��ܴi��� �$�`�#3V{�'������zY�[X^3��?�3��^Lp��~g�����-
N|�K.9��j���Ή`i'e�m܆W$#+���c����zq�- 2?t*��������-\�rL'ߺ�U�咦_�����!��:�^����
1�p�Q2�}*jרq:�AA��ۚSzF��4����tT�5�C����˸,,���ko/TɌ?���!P]���tQ������V�ig���9K��oNtê�	���8�^Xc�^������҉�;�N��\�HZ���	�{m8��췱���-3����� �� ac�&KI��<#^Ln��|���&��s�@'GvMlr�cʲn�� P	��~.�\��?�߂�����ĵ�yO��>��)�S+�z:X��i�6J�F&˚�����f2.ٷ4OC���f�p0��?a�\��K=LU@T^I7�"j ����ǆg�O�u��
�����c��\C�_���n��)Z���}\!ER�P\�">D�L�p�+��\�zVÖ��a��AD���6>���y���!E����icV��ABv��:�N�#�{k��f~֚��H���-�&)� ?,~��H1MԠ�/��/n*3�G��?[��!D��5�	'��+����-��� ���c�8`��۰q��[�>4O�'�_1m6 ��e�ϓ�bx�X�&b{#��I�kf������%e�K���"l�G��	 ��N.�r�VA�`�u��#�Ѥaz�@���҅$���m�J�9jpE?]l�F7G~ʐb���]�3�A���k����yi��������/ǩFE8��ء�U4�5׈�������`� ��1�3��C� е$�|��H�J�v?"f�4:ᎿϐKɛt��8��6d�2��j�� |[ƭ�
�bR���I(
z3�n��^�H7s�ԉ�����V�*��TU��5ԭ�38*<��Fx��,����-�.Ytq��ۏ�4:�F���"�ۤ��� (��U 2�̋�i�V,�pI�OAѦ��	ez!ILOqZ�d��V�"]Y���W��v�7�4�{�+���8�"�k&ـ���K�K��g����w�\�l�O������V����`�b�HB j��i~��ݡ���;��0y��Zv�"RhM{
OJ���PM�6|�;���G!�!��S���˟�7썘M�eY׆EЖ7�t��v�2GIgB�%���A��΋���b4�ૈ���/i8�z戓����Hť���ϏS�X=��"��
����Qv$T�LR�(�22b��/_��&7�Tp�ʁ	BMb���os�#��;�8����?@!aT��.���A��f�AgTG���Ƕc�Lh%�i=Y�Z�b��G��)���:~�3R4��2���}���3�9c����=P�������������xp����S��a��v��A!&QUD��%R�EMx����ɋ�]��F��VH�Oac|����2ɷ�~��M�ԀN�r?����e�H�$^J��c�=5��������r5uo�K$$�P��b2�ϲ^+)��RpVBy��VV�H4@!0xw��F�-z'��{����75�X_�?�װ�S��4���s�۳�r� �^ʚKe�^���d^�UWX���mP�Y���0���v�~�)�u-1 �e8�����P�Fr]0��ĩIT.SX�I۝�� z�[�m��X%������4C�IՏ��ʸR�K�4�s��J�ĦA�Ӫ�]2���V�f�0���\�M�d�g���M���R&��Hj�bF쩂��v%��HK��?����	�N���^�z��2jcbV1d��v˻�6�{"����(
nb��aw�C^�νd@y5�K�$JX$�3�7/����Џ� �M��f��yMs�v�[</0&T�r^h:9����� �w� ���+;	Y^8oj��� ]n�����v��>;O�iP�$D8��WJ��K�)}}3���ou�8������hF�Ƒ�b~8�H�a�fg?��B�3�tkC'�DY��!VT�0G�ݴ�s�(u��{�=��"�ww<I@_˂j=�S�S.F˗�p>Ӂ��?��=7[DžI�V��z���;!*�+Kl����<9�ԥ���B�}�P���`��om_����~������|m�µ�@d�,Bw��8WB$�d��<�k�5�@���0����Fyohy���)(�eJg��Ns�w�N���f�`��Q�lH?����&+��)8I@\�@�������.�4��O�w�Ȇ�)�G��b�qI� ʨ��ep��/�=Sڟ��yK�P�uٝ���]X���!:�L�d��-�9���@V��(1~"� ��!Ӎ����Gf�'�E�*��vp�$�U�xb�Դf�c|�N�@&VRWs�xkrU��S}����U���v�N2�������N�Ր�^���Ҟ�n�a�J���
NAk����sP�t��F�{":	�L4�s�MQ�H���r!BD:�^�{�f�S[h,\Yi�� �-��N����G<�JU��w���;���Rϙ�ɇOP��6�,8�s1��O�OB^�Ԍ�}g�Y�X��8�c5VeO�.A��A?�L��iZ*��U�U[�N���Y�5�,�v��|2�I�gވ�͸�2A�E�_��-e �/�&�0}��;>+/O���ȵj��&���W��"��³�9�����?�z(�<pD����=�����7?J��� 4v�Yz�b�$)�4&�W�����C"�0`z�=`v~�%b�jǚT�u��P�Ɛ�k�'�#8�2,�nĈ�eI�B�κ�� ���XTQ®�`*��#��kzx�8�������=�������R�t-�,7�J�� ��Dě�b.����
��_8y�0n������;zZ��`�މ������� wEG�d���'T�,w@�b���v:�c��H�ۺ*��ѷ7����X�ztF("5�����y�rS�n3o i8�<���XgT�%��c�
h�~Z�%����j"W؅�uO��HR����A@%�>�q�zڇj��+�<����� '�\���ۯ7��qu<�٣*l�6��8+6	��!��=�Fг�㦜62(�Z��˽����?u����bإ�2�(|/H��A��@p�����4k��5�4����d����j��� �S�J5�!?��ג��Q���<��J�!&���Њ�d�6�c�gy��6<�JDJ����YC˷�"����ۤ�V���3�mU?�ӭ��|�\Ѭ���tk ��CǑWb4BMy�"5�0�����z�.+�6�?����*�HP^2O�p9+��ppź3(p�(%ο|(gE���؃g{zu��B�N��a�9�_������@ʐ����/qne��.���D�L����l/]�fg�H�'����LmJ�Yy��S8 �Q\��!��HC0�u ~�]�EEQ+[H����o����L�#�K�&I�C&S+a�̻X��[R��Vl��4����x�FKhӮ98���,եϢQ� �7w�[�d�_���m�G�Z�[N	�4(r~];��R���^o��&�\U���M��U|/�#�(@7z�`�Ҵ���	��4�c��%w�⼝MN��=�3}�
C�k��65i�΂�óp��4#xZ�a�o�:G��,�
�x�!�@��S��	B����JcJpTeG�Ҫ���	5����|](��p�pȑ������$}*�ua�t���w7d�76V{pRIB�����xTn��I�?��� ۑ��n�DC��o9�҉�9>��/A��փ4�<{��qt�2��x���Z՝t%!����ו�/����Uw���>�Pn�?_�-R<�nX����������8h���	�"���`�'
��; �V���_��uތC�z�Ⱦ�xNd��)�L~��φM`_i���[1�Bz;+�u:P����m\7���aӰ��D�)�Au���f�ԗ��y[�Ŭ肬V��*G�[oy�F֓�x��`�ꚹ�HA�� ���*^g��"8�B�8#~t���6���8[��KR������;&m?��2tYZѸ(��;~B�9UVM0 8~y�R���m�m�XK�E�L��-�7�sB�I�|x��y}!��/�̪�n���](��'�8���u�P1���ƨM2�s�.�dL-�2,�HB7�'K�\�Ɣ���u�\��*�I�����t�����s� ��^��W���(u\��OUI��#+��*�.�*�K�}(Lb���/.�x���ވ�j���2��R8�&� ���d���.Ä�򥥏���Mɀt1�Q��1-��d/9� c�dƒ$$���1���v��Y�q7~�o)kƃ������;���h�!�_RP$��" ��w�ߠ�"M��p��.ıx��6Z�;2qf�Yp��;VH�zE%r�3�T��Z�����05waR*�
$��O�m_YAq���M��j��5�cZ���&�ŵ{���«�n�3to=F;����8�g1!f��$�_�9L�����0D�.�{�?y����� �i�gj�sej%4j�3f�s�.ՠ�����But_'I>�"`���-��,I�);�x�,jI�wn&�,q��љV��?���N�D�1���C��k1{�Ŕ������D��vu�於ᘃ�Y�^�}����7b��C�H�,��;��s�\������`�T�se8���<�6B��q@��0�,���Y�W8ӹцm�y`��9�#�-x7We�]*�I(d.���� ��XG�B�>��~�+p��_Q�G	E+.鐁���� >��>)�\������!&,釄�����HR�);=�P�z�5kO�	���H!F�|j�����QRi-�O�����RF�S��Y�M�T��/�q\%�B��7�f������-����R=��YW]%�~Ҡjv�.?�}u�����b{~�.����!9�du-�� �|���p�x�bܦ1��9���\Щ���sŴ`�(�wŲp�ɏN�.���Ų�J��p����G�r���[G�<=��
�W���wv-�OEÐ	Y@w,�ILW�Z�
���㜷���z��d�ݡ���r8̍,z�M�p�.Ąo��߼��8U��懩h�r�Tfu��s^�1s�m�"	�Sų��o M:�*X���ժEN��'ǫ�gֶ��� ����Ԕf�������"KD��<����W����q��'0��[s��֚O�:f����K��8����xd�A=ػ<�`�BX,ʒm����A��愸��ƥjNuN�ԝ����pG�$�󇙷��f?��0؍D	�g�i�Fwt����5t{	C�`���܌�F(��p����\�aX	k���$�O�Bf�Zۂ�?�q��GܟF���.�IԈ��0'?+i4�;��"�R^�0z�� P����D�Nh_������tw�1���9_���'x;ؼ�ф'�v��8p-��֖�~� M�j�g�ſ�yO="�yv#K�{kb�&�"�@��}����l�,c!�m�$�+t�ٚ��=tk��y[�=�x'���}�ޗ'?��t�Bb�-�u�{/j���pRh�72��O��V�Q�ÉK| ���?��P_^S!��|����?����5vo_|���a��t���4��H5�@�z����5��8}��߀�-���$lA�ަmol��C&�@�9��ox���"	!�fg��wg{��}�j���ԉc��"L�����:��䪃y����rM�����		K���|�T+
Z^�5O�𜗈.���PB�r\�j\�CۣE�H7+]�ב���&�=P�N)����ݎ��;cd5���7E	���Is2��*�L���f�-N���c�Qd����t,;_Ƞ=ԣ�7񜊍܎J*��5����&�Q�������7U�n2/��(�y�*dȖ��6UP0z��$��c�P���
֍�Q"k_�p�fA/�)7D
=u�H��͐���m��fV�%��ĜǝVp��`$����[��`c_<!������/̔��7�8��U��.��6�^�CA�k}a#-��^�`����d&"�g�W ��_N�![m��3'�g�G��y�š�B�&�dlU�P̬/�\b�����t�HvOR���[����Z#sPW)�77�7������j[���}��l��o��fV�dC<�5cR�Qg��ew�W����65�����lQ�\�%a׍�VcSI�����H&r�������7�45�L�'V��X���t�mr�@�#Cm<�{�[�ً%��SS���/��ʓ���xg��DgL�_s*P��Y�k÷�ކ)9�U1I-�!J'���D�ܔ/d�Х,����O��R\�v ��/7����z�@c��$.�;�}o�^^����*f�g����X���Jg,}�G���0 U[��\:GgA��(Ƒ��6�#䪇!����H$˜���y�98�ƁI������ךฝr��z�Ui��NM	��l��䒛�1[�\�;/[�k�����f��KȐ���
M����J�g0b�W�\eL���){�m�37Q�'�3M�
�;٩u��-�|�_u(�G��G�������V�������,� acF�����T^���(]5�@!:$،-k����V���Ќk�a�۹ZfS���,��] �G�8߃"1|�k!�	^��dk�;��L8�����"J�y=�o�-��!���Q9�g[�0���8s�$�f�����ԧ��1Djf�>��B��Chjj_�`�z��&U&a*�R^A�n;�]��Ql�.�2ACS]���	�0�(�=i�<v����c�"4�����3l��+�����?�0���b�4V������H��bX�B�����n-�D�P�z׎˝/�6��6"�z�&04y0,��G���wxp�����x�����s�Ơt�C�?n��I�)R.�0�0u���ڔmʈ(�7��ؓ�K$p2���a���������h_���E�\瀲��&��A�nh%�;1QRr�+ǹo��D�jF,���1O�[��7fN���p0���Q��u����/*��pq��g�e�N�&J�$@!.���$��yN2���{�z	��p�O��Q�Ƞ 4%[1���8�o�bXR��S oM�*z��nU�����D����G�b����裰� �O�g�\�����c�xqZ���3��m�;<���m�b��y��3O�r8���5G>0�_�)��0EY���#��+�t�ο������S ���2�%H=۫v�K~F�3I��,!❌�����;�����cLsD���J��d�z=V�M�|�
�K�$��\��,�= H]��J�;�/mႾܗ�c_�B0;�V�}|��,/�8T]��9��a}�X�Xؠg��z��fh�����{�dǡj�? T�%��7N|O6/����5��Swt|W�����v�de!���m��r��!�R�TQ���É̝_����������׿��)��r�	��y�,��ۨ����~k����PT������ ^܈�d�+	���v19�b����R�ò�����Uf�|����H/z^�K��w��B�����Q�>dY�i�\�����R��sk������=u�i���h�<��2���d����jqly$��=�#Hl �_��]���ݣ�1�.c����o�&bڞ���7R[�!��{Eq�ם~���~�]�<R�X�_�\�;���E+���L�%|MNq�Q��}�wnq���|��RfF���I0!�$@6e�Y\����[ V��2�c��J=N�vF��N'x5�#@��Y֗����V������ ��X����}�x�*�$r�b�pC8��Q,[��*����\��u3����'6Q�4z;L`���:E�sf�#�KA:>����y���a������TW #��$ t\����I�Ӯ�yz�fz�����hq�6	����P�`[U�����,��x4��D �?]%l�<%d&�T��M�r��C��:���
���)��!��=v�剂�WC{(ΐS�N}�����!!n	;���6�f�[��fCzа�Ja!n�(�y�|�͇%Z��UQW�~�һS��b0gB����������N�@,	�а��z`���.�A8�4V <�sj� ������x�ٜh��jUnh���y7�$,\,B��:���C۵v�5e�q��'0p�֦���@���Ϩj�>dԧ��$��;�0y����}Ain��G���2'���F׳hO��I���"���T\g��Iκ͖u@�F�������U�E��s�
��;�������}�Lү���B�jĨ�J���-V��l'"P}Na�mp
d���C���:ҭ�8�X5�lX��%CML���(~K��LȨ&K&����������s4���6�#��V��K�^r��}#����;�P��X�N\D��o��u��l{��AIQuiS쟞e��Ѹ܋�I?�T���m�N�4ã�G�l:w��`��zE]<�=ᠩQ؜�i��6�Po��J��a�=�yP9����ώ޴S�&�^D+��+J����TJQo!�;<[R3�ƃ���&�}�7�R�@f��A;�sTCڵ�䱆�ZJ��i�U�g��&NYٹ��F��9URY��zx�������0j{0$O\#�+��t�3r%h�-�^Uh�u��p�t`C��,H|5&g�B�3kصM�'K�mA���gcG��\�hȌ�=X�m��������P�*��y���S�:��m�H���7?"'��=P?/ 7�m����Rk8x��ous�R���7<�k��5�l5 �����h�J�I���B�<q� �~<gT�˯�y��1������	t��9�����24Q2�\�b/E7l2@��� �+u{w�{3Ǡ�'�� s���{��񦙈4��W�o�e�� ���geL`@R�� ���1s�����.����hl'�cQ���5rb�@����Ԙ��T���(a�f�S��Y�ľ#��` �{[�v�P��0��GdD��f�����
uUӵ�څkF�i�O(� �v���m�>Z)�Kgà�VC��X��2�;H���,Vx�@�)��h���C��� g5ݏ��Q������V(QAI"+��@Q�q��^P�ΦQw|�Y�'g7�r�%&��Y�d/�~���܎�ϡ�a	1إ����U��]��}�}�(9�r���b �"�� p��X����Ԕ��c���6y�w�@��t�:��o//�&!3�|����P��s �U� f�1G*�JJ�v��zS�R�э-Z�)����me��JX��D��B����6�`E{��8]��|�*���[�����1���� /��u�많7�����3>��``�����V�_��t�˾��I�����ò�f!9ly��]�3�m	�k��2w��[^5�2$@((������?j��Д9���˻�y�z�ܡN�v�*��g=;pdv`O�/`��L�����0a2LU������I=ä�Fو(Q@��{ �>a\;�y "Rx����V����,���Er�;���S��KlWC<_�M��� 30��y��n��E(Ёx�=�"�_#�/؅1�����0V2�4��$4�Fg���qو�w��[�����f#/��t��.U��Y�WJ�b?�2";Ɔ�fE"��vX�3���d��"���Ed�0������N��S���c���J35o�N�g����m<<�^i�c�=yMT�O�%=L}�����~�یDY/y}zc
�-y��_H2�_!F�O�K�Q���|���@A���ه��Z��\�:�H88�/��6NꉸA�fp"����"��9'�r�w�	1��_#�z���A����1bm��"��������'�C��>=�~׫��j	α|��x��?cW~�g���G�JN�� �ׅ�̰��t�gy������.MۻʰOz���Ek�0� ��A�t�ߜ0����ÌJ|Y�69' 7T�у�c�s<�X�7�[]��.
NO;񵺲!0���W�t����g�~st���0��&�oיUi�7iXK�W'WC�,�T���q��0AU�����O�6ǟ�J���b���94.�����)��hu��a��ȿ��-83�i�>�O ��:s�
	�����{�ڪ�������� e�k��&K����a�ʸ �n�,��`��u5�	V?�ņ�tH��/��9�=3�R#�q��9�x$t��1�q�]y:�ՙ�;�.uA��z���S��u��QV�.�ѠSV�Ù_�y��t@�&�AΝL�WT'&�C <i�����VYP���a��J���p��(6n;F��f��q�&:���_�i����UGٕ�=���G�� b�-��:�i<�M���*<��Y�R�97��	�¾S�=�9w̯ˁ����Tu�t�5h؂"\A���7�t�����b��G�P�$��Yp���&8��y���&�������q0�(��w����1�� �DX:���2���T}�]D 6��^�):��1�Htf��vʘ��ǝ��C%m���*;^E����(�-4��Z��k|x	�7yt�I�#a��)�*+Z������+��|�/����F`���P5o:z��
E�N�ɠ	-c��{*'�r&m�0�,l��h�o�X�9���7��;n|~��{���P;���q:�^�r�B.��ԮC��:��'��_pDr	:z��*x`oG����>}0S�ԶWwM�6���u��#?˦�0�X�I⻭�"ο���~>�-��	�0ч�)-J�2�[���) �X�e=�j�{D@+�M�O,���>��Ԉ�oī ]#O�|]!���Ig	-ܻ��V�ղ5�ZQYig�*@�?�|������{�}uU@ �ڜc���d.G�H.���Φ
���˥��<,"#�!{ċٷ�89Ř�c�ip:��10��yED:K/@�6@�ȁ�%e7�1�����d0UI�u�m��u�C5vbF,T��0$m�ī�2���d5��{�l]x/W"��8x�n��d���6���'�p��উG':�U6��foǻ����xD�]����@��W�<�,�c%��&���k}q��Yajş
��7�j�<�'���zX8׿0^�B��*2����t Ƚ��q�̫処,��ُ�W"��KZؠsl��`��J��*\�_���k�+��Gqv�
��-;��g�X��L�pU��X�(@R�?�3���y�`�# �����&���躀���ܮ
L�/����%��)e{���b���h݊��w�/2i��	n�9�L"��f��~1�&Õ97.|�H���L�� i��iK��ie��,��q��y�;�8]@QpD�9����5�j��&��<:�|L�RW�<$�Z�|� �mt/=��؜����w}�����9  г��*Y�S+	�[p8?�U�����\���*��g�'dà�z��Ub3����{��rU��{��%��1�Q�EшV��mC�x�6Y�)�s
E/�*<s�9�"��%[�:���?����,��s���F�6�e2#�crq��S���`�7r���φ��ha/z�֩/���H�I8�8z��?�J���8���/ǻ��IJ�����tˇ΁��e��o�T}���6��{N^&#��jRO�������=kwm {�4?���uF�>��9o����#��Nt��l-�s����n@������bа78�������"g
�Nu!��9�7gS��Pv�����f���VB(�*����v����Q������28���vU$��DU�F�Ə!��D{G7�!�P�M���&~���SMd�	T;T%Tc���׹�vZ/M�b=�R},yU�!��-NeҶ�L_�l �y�ء��o�=��K�l����j���k���D�+�N��j%	zQ�ڏW��}�A�~�QƵXp��MGYC��?�C�z�g��he��$��]f�}]�.��&�h�I��ٙy�j�A{!�n:uTrV�M�4�E�3�8�Ur��m:��uė�(ܖ2��Kn�w��,p���e�#�%۵�OU��<y\��k��Y������2��aU��(4�Y3�
�k�1��j7q��������3������x������v�X:���;�W���_�e���uEk��9�1d�A�EYJQ��`#�)Ș����w@~�߁�e�_夊�ƚH�9ƹ�ڸ'�B�������1 Y�4U�8�cM��6���bn�(���V9��6 @#��=�HO���b#M�xj��AJ\�ä���W��J����@�d���=$�0�DYU̍1O"ei��{4���Q��U�o�$7U�T4[�	Z���"&s���h�&�w�ۛ�	��o��?QW�=��,��{�V'�g�M,�bՀdR@u�"Z1�Nȸ�LA������#�TS[����ʘ�K;��q��Gǁ��b������"l%�����p����Rmp[,O^'+܊��̕��eg�n��q�b����U��":! o�z�ޥ 4z�ݤk����N�bY�#������Y�
W�+nD��u�O�"Gvq<C]�(�s�x���/OBۘ2�[�0>%e����Şx�9�w�-�&:��q�������y30h��z�y��*�5D��Ds�MG�"ğ����;��/�j����́A���W��Y�ʛ���m����hՄd�L�Rez�<��6��I���'F�����,t_/�J�W%�S@���?:��ب&(
s� ��A�����Ʋ�=�1��qIfEl�������W��Mȏn����"QN�u���]ft� d�3�~$�����m��zF-�q̣�<���"�Z;��zk�ñ E~ ����ۨ	`]�ͭ���Xv�9��Y�(2���^���̡��RM��D�f�G����Z����O<>!{Ͽ-V�~snv�*�)�R��yv0ΒsָYp�@��Б�;`�Uk�S�w���k��6��2S��Ԩ�'������V��'x�7�{lC���%�n/r�2�P����}\"��
5bs�=wR�q:����.����;�d��_����DR󳄎���7��/�A��Y�A��U��3:F ӓmK���v�Ŋ|�cI���vRo���ǳ�rH{pb�RB`E�(����%��yF��������md3 3�U�WMn���� 8��� ��h]L����O��1�+ú�m`�f��u���".Ú-�qnz]K��lF�;��������_w�E�A��7E+�N�@��֍��!{��+\�;������&�9W���{d���'��7�L��{m�c�R����Iaˡ3������o�V%nؖ��[@SCAi�\g���	-�d����w�:�������r��܁��Y�6Tlm2J=i��$�������L8��kp�! ��Ǧ���}Jv�ȱ�Ҳ�!2٥5�1P����� *��H��5���߰G
̈́,�ќnD�E8XJvO�z����|SA�(9���-�������HTz;ߒ��K&	��V"F��̩@�b&�`�bآme� '6ZR�\]ݲ]�Ģ��}��c��^u[xY,��	��W#���[�|]��o���1��HΪn�bsI$A�D�
�`CH�������>&ʇ$�$m���ؾ<���g����i�"������K!Ư\zr1�X��N���Z�P�������Y��bl/�|����[%
�o�=u��������v�
�.����ѹD�j;s�YN״̶�E#��#���JQ��S�7��%�bk�s���y�v.P��6HG��e 45GQ(�k��I��7_��h���r���Ib��⨡��p���x:hc�c��Y��(#��Ɔː���sV�+����vec})���yG4_~�;=���ˤN��U,Z'2��A��\^����v����n,x���1��P���B���8�I�"*�E Edv�O����{g�e�Y�b+�(YP݄�;qwV�r�s�(�C�8��m�G���ވ	�/(�z�v��ᗼ�(�������߁5^����t57��e��i���W�+f$a�;b��r�&!�!�c�m�¢B�~#��zBN��>l����K�D�5�0ԓ�I��m�6�v���fX@߳@k�k���x.������3���뷽����lW3b[����k������2��Zu����oC���OC׈ '=���K���b8���ȸ�N��&����3X����c�
&��T(�f���.����	�
����r�Jğns&�E��<g�(62���Il���@�cG�;�E��8�����
���fW{��J�˟dv��j������S!��Ǟ�XJL�:�#���[�~E�Iw�n:bXԣxP������A��Ĕ��=�8�B?P����O��r4�Q��61'�B;^��}^�`U�a�θKg�ץ鲧�W�+Đ�8.�2���~INo��Ķ�1���~/�� �A1�f��7��^s�n���7�{}01��
n�-~�bjל˜���Od�̰?t��0T����4�P�g@y��e��W�`�q�t`�څ^�Ya"蜔o����	�]��L���#�3��r�a1j?��u0�=[ڗ�{v/�>:>�� ��!���+��T������u^a�\o.j=�*�Z~�e������|ݏg�b&4����Ys��;���jn�}Ҫ���ڂӈh4r��y*���:`�x ��'��x�`���,K��A�i�l�����<~���>��. �����U	|�֛YI!��������B
��*X�@�E�+�w�����}@�v���G@�l�~������z^"(ǩ���	1%����Dt^��}���M=���Y����@Z>�/���'��dvR�뒭{O�6 �����&�Qcu$]�����N-����<	������r���[��(P�H����Er��9�e�k�(k�xڑ�m!�Y
�^'Qs�>G�4�8�hy�B�����ŕ��+���ͪ�H��)49����liSM�9;��©�%T���F���Z���0���ig���r�i�&��H!@X�/�O��NV�d��=�G$[q��x(��k��
�+$�G�O05|X�3����o! q�v��0-�),���������Խ>�CZ�%J+1���� ��F��9g��r��ӁK��1��e)<e�zO����_��
!hg���܌�d��Q���~{��F#�zfM� -=����So7A�^]�"��s��2�5	���:׭&x��<P�m�)O�rrܠۓt�?]��FǺ��3�=�3��t%�T�i4 �z�j�jOq,�j��V�Vѐo�ڧdֿ��R���Ŵ��ឹ�Y�}�ߚ7e�����Hi��]�i�gmF���l/O���y����N�rP�z�]��%a|l�?��˟v٬�����9|ĸ��,Ĩ����p����2�1�oe�!3v�jOo��hp�;�]II'���T{Ps�|n�9Bw?��n�F�����~<��/{�<7�+&�/ف47>�d�omM�������2ܯ��I��}�C�+�ɶ�χg�"U�,�0�~!!���;��5&�m%z�y*`l�h���jD�Z�e���c���:�PÓ���m���q��j� ��\�����}p��KW��=b#��^[�x�G�4�i�m���O�!+�'�u1�C����Wa��PQVL�+�y��4�$�����]��򻍟�ȣ��/S����"^Qv!懬�(��r׫t�"�M��4���\��,[&�C<�_Rı�$\��Gkhڏ������K�\��l�!��i��!g��k�^��}c��?���z�g����.$�.��o��/��^�R1����~ݚ.������{�����'�l�͇-�6���!�`DA)$[�2�߂��c�}A��Z� ��E�.�NC�[a9�eq��3�����=
���t�ة �_=k��.PE�fQ��S��<���e]�p�{�Z�y����h�9GOڀ�'��h�VArF��������"ɸ =#o�a3����O��dH=�=�mt��� �<i�6�"�%���]�$HUF*�6�"��lo[]��]�߼[l�+pR�Ű�S��9��&�������]R7{�X�ċAc�3,9��0��]��;rБ��������ǀqC��Szd�輠���s��%BMx�SWa;Cp��)�����a{��J�.��M �T�J�[���&}�����'�Ԑ�9�����_�uA���g��D=P�OV� ���-�:���[@��>��0|k3�DT(�潰����CS�޶ t�yh�|���|/�9H��0��
$u��O,K�mGd�X�No2ɪgC)� 	?� D�[��R˾O�TD�o��Y�	赪��һ+]ۻ����M��,r��|o���A������@6i��8	m����b(�F�N�<��}m����W�="�8�^����a��ۊԇ�銭� �p��-�)u?Cpp�ʶ�V	cគ�#+gn`ބ_�in������22b��'� �d�6�6H[�0˪F���n7�~�	��a`�HX�=�Q\���z!�Ld���MM�P9}*\zΤ������[�i�����{��X�NXu�NЕ�N�5��&$B*�X�~,�]�T�K���WZ�����V�h�(��p������'�,@YG=uouR<�|q;_+��K|�ǀ]���;[eAђ�k��a&ܗ��5�gS\2��]ͩ������<`/p��劧����Ev����'��y���l
!���>��U��I�����sO�� �ک��Q�^�Gۘ�&WB���C�w��V$c2]�Շ�_#��،�F�����M{$Mz�xwkC�M���e�̫�'|#qN��\�g�C�[�D�9Ի=�BD�>{�?��|�q��QЈ�[��4��C�����JWa�6-�/�¥�����I|�MQ���ra��h/�YP�}�,�M��AxWo���c��J��qe��*�P���t�4��]D�xA�]�n��&V��3�V���_���X���Ap9���:Qߌ�"uP�Ɛ��_�J�iX/:.*�A-�����<���������)9n�?:�j�^�	�e�~��{8'XZ�f�&4v)���]-O]�O0p�܃����t���H�"{ %�][��m^K���[�" G>+��jѳ��"��#ߙ	�*BIXqk�p�q��[صM�!֑$ސs�w����q7&�p�1���J�F�A~� �&\��C\L��ˏFRb���Xr����c�/B7+���3��{��	u��=y��K��oZTf�-P��/5�+�2��+��ݒ�3ڮ��!��<r��{�AP��|�퇋.=Y£&c�]�~>��6�T�*�>H����z���n�P�n�FBcG*~N�!��K���aߧq�3f�ҧ��*���w�����I���&K�G�a�4�I�-��$���t6���\-�|\V����DH^�Ju\򕣬�A^%�
���7'"�y�_��D-�A#>�֫Fg���� mF�ȱ�>?�?��C^�J�CC�Iw��@��;~X���}U���?�)D�,��
���W�'�9�\�SM ��o�&25�!:/�vĻ`=_@�k�6
P�o�����o�����^�L��[���@��mn�g�{�����H����pG4��jwS��YZ���2�3����3X&�D�o����%P�˔�E\D?e!���LP��X<��
�/��;�i3�µ9 y�W%]�fz}��t*h̫⯃	�at��2F�w:��P�%���3��C��]�����9��هR��wg�0%��l<���LBDQq8llSo����٠,�Z_�ӏc23��?5O Y�fl@�,�rD�����F/��Z�	II�7
ȩ�$�� R���1�ºo%�t�.4a��e�v�����zc�x]�^�+�h %O����������{��jUbO�
@}g#�{h�GdVa�q<��<���&A6r�O����^�KG��’��� ZG��l��qR#�tsPEj��Y9`+m�+TsE��]��u�D�}n�0YP�v&0��&��4��	Ŭ;���s����kw�µ{3S�l�M����X��Ph��z�j��i"�5	����N���i>�嬙񔲤;Qu�~���m!WX�-Y_	��reW~��~$��R�V��3�׷?�fu�|��H���3ĺʊ�ڿ��:z}��ڸQS�3���R�����W����Nss��^�E���C�c�k���7��5���-��O��
B�浴F����d�;g�3܉AeFk�������!�Є��̚7����f�jIDR1}o���Um�����T���Ώ���Mq���𩇡"��15�?��	j>���� ���C���䩱#�
(�l��ެ4O�*֎Y��c�[�8���L����Y����U)��蘂��m�ڎ}N���S��S�6ͺl!w�#?�@Μ쌺˚�`^LP��]���Z�W6x��9�T���bȚ*3U��+-X�߻CLY�ÑUw�1H&l���� ��Jpv��9�d��1�·2��ˆ�{/� 0���ʓo�\J���zƔO\3�"j
��~lt���V2p!�RF�ضM��z���iŸT����ѡ[[��_����w����7	���O�|���W��V�S���D0��c՛����Ȇ���Jק��,��9i2�-]J����/9)�KNҬ"'��Q��G���W�_8�SR��w�X\���v!�K
��Sr)ʛ�ŵ���x�O`S�F����ٻ��*b���~��)x��3��tFUS�az�l�wZZ�N��tCmS��A���jN:�����������d�}O�p�6���J@�ˋh�ԫ�Q�b
Q>R�j��9�r��9�"�"1	��5:�����ԡ�<.:
8�]�w���"�J�n�X
M4K��_l~��K.#<�MCJpR�y8�/hY2ܪ�iU��߿W��7�S��Qm�x�; 鲿p�p�e�h �@����kE��XC�%=��IB�IzE�j�-��-�Ky��:8c��aPTv%�\����*ե�u�{����@�P�f1���a,�l�([��u�w���)>�ż���a��r�o�ƚ�A��$I	9{��I��b��u��-���uc*�s4ӛ1�Y�}���lN�n=�:�X$�e7,�$53LV2�h퉨�7��7Г�y �f:>�wD��I��
���a��
��^N��H�
S��^E���g0�h�X���=�_{���[/���{��}��{o.f���s��#��>xe�$�E�7FZAj�aVg��^�o������ǵyFT^ީ���,v�,��wt~�j��V���Z>�A���2H����O����> =�[f�XTy�E���q���uO۶���G0m�l�Z�*��ыt�=o%�'ل�g7h�̯��n�ևz�:�R�Z�H�2�.=(%�;�\��7S2Iax����ǀ���u���n��SdO����
V,G���4r�oq���Ϗ(�ME<��rSJe�	G���&��03��B���=�����^(���S�4X�q�z\0�aa[ +�G��d���`x�C	U�ts��M�B�d��=.�tu�|���I�{����>�v&,:FkPk��ɸG�9�*����#_e0�ϥ�&C��\>]g!���ɳ���>zy���(�{Y~�"�ߣJ�������XT���G�	�3�x��I_u�m���F-r"2ؒ�ʺ�ƺ�
���Cߜ�R��'e���p-�涘�<i��׽�ī��}.�i�wE��1 w�k8HH��xGV�5�P���J�I�|��%�,I�gP/@�#3P^./W�'���u�.��^�w��4-=F:h0R�;9��Z�%��h��'>=�8�*:��`H��}�iX�X�����:̆�/�d�h;Ls&H#o�� 0ͅQ���Y����L��v2��f�F��"�DI���]J$����0�ߣͭEd���/[�I� ]�	�#$lP�JeL_T-��[)B��}Q�3lF��@��f]�֥̌ܽ5�1H����-T7��M�?�m�>nuy ɍjF���{F�c#<A$�>�E��!���3<I��Rm�l���=hۂҐ���G�)���\�Tn� ܰ!�%�̭Z��_^Y<��qݯn$U�q�ܰ!:^7��k�7O �*�LN�um���刣,f�6��K��3�U����3�$�V]n_��������|� ���)�E��V�e������4���c���}���n;߇��U�4nV�^���[0����]ɻ~�Q�9�]2; |�.ՅU֕,@/sU Ut�9QNl8F�d��Vc��O A0 ��q�R#�]��ՄG�y��i�i���|Y��
�ܖF��u�   d��y��_'�"c6c2a��n;�o�<~l����J�w�;������b�p)��	�.����!"��ώ
֖�nÃ����`k�8+(1�o�ՃК�E
~H�b�J�����!���ޓc����.�����R˯����� ��|����N�/�q�1���I4���ޟ�Y˞T�e�M��$�Fꏃ�C�/.`>@����qU�+��ܧ�W������ӇQuPB�Z�)}�d���a�nݐ�ɘ�������L��r]�`ѹ�����a�9r�n,�M��Atf^��5����T?��^���;_~|�E����v�\�gB<n�r�京A��s{�xA���C���W���5 j�=�dXM�5
.b�!�����<Q�lCƈ�T�C^s��/�T�
���7�>/�����H��f����N
Rϻ^�8� cuL:﨣b{U�U��}����8��*x5ϵ/��O�R�M=��)#�W�#"2�G(_.�����&���5(@7�yU���#���^=c�O���%�}��M\ܶg��
���IR[��5��bț�� ���1�����:��I�M)6�5��l�y�!o0�~�2z*��&�se@�&&S��0�7-㷰��1.���pn�l��:�k���6�-0��h�+����D[M������r7܁CbxKf����E����+��|Q~?�y�l���8�`�Q��'^f}��u�cҨ��q�`�4%@lM�>����ȋr��F��^}v��;�3kf�г<:��À��-��)�]@^f�t	�0s&��
��ƃ�����Ξ� Q�#��jPD��0����Z��b7��&r�_���{�)ٚ���m涽m��";�S18 ��,�'�O���z�W#�G̽��Tn���0�h�+��H�)�Rj��wG���jiA������>l��RDJep�#�0/����k��C�N2���n96�Z�'6�6���d%�����)��M~�Q F�
A	Q����e��) 3�H@O��������z��B��/��.u3͔�ɂwb��6��_�a˃؈�xY�R�f�:�Q�����c�{���_�~i��#JF,/��!����7��ѬQыB9E-�vO�Y�ϻ%*�O�vPK�Of;F��T�h׽l�ύ