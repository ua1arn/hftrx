��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ���7�dA=��p�Ȥw썀S����?8g�*��'G�>�����=�1>�b�1z�v�'y��)��{�2.��R_��]JLJ�D/|왒^�V�u�B�Qp9[^6}�	��7����M������g�]��F����%(�ȃ�H����y���A����PP0��D9E�Z����͠����ye�T��~��H�e���߫^�d��z������4֙����̟�uk[+����4$p�%����K�l�V�ټ�[&랑�FN���Tߘ��:�UшbQ�f�����~�e�B�`HH1`�0���=#�F���n!�L
}d���\�2��H|@��
,�Z�_���t�����B!��S��
}����w5�+)� oI?`�WW-�W_��g���E2|\Qj%+������Ng��%0z ��״{���˹У�+��D>R�G�}F:�b�Q�)�M�N������~���(:o��3����Kb����
�h_M[�f��Q�Ԍ�05n��H+$��sp�-�ЄI��D�Gt�G&�~G��"c�k\ �Ck�%rh�U��M��|4����zVI��aE�ާ�3�x���Gx�h)X-YC-������^�~/QP}��Vv���x�I�i�n�U�q��<L��,儻!�g��mYYS��ӈί��=2
a=�ӡ{��&�%r>���A��u�,�:Pzo��=��G;ړ�y&����Re�zR��=5��A�����)p���Br�gV��n� �oy���V@S o#�E���t�����^�x
��M+] �E����Y#k�f-�2?u�#�~�:7y������?͞��m��jӣ�-�7���]�Ů%{G��Y�n��X��½�)�b�UI Kvjc�l /Fg9I�r�/g�;��LJ��D)�;��.H+i�˧IB����:c�OG����\!�"!q���9X�fv~�7j49�������^m���KPM&&�c홎]I��5��د#�F;|�s��A�P�#I��w�P'����V��DCO�����>�������"��&=h�.s,�?19d�����E ����~��VZ���e��= �ܻh�b�qG/���g,6�q�p�ٜ.�&�u�ߧ5o������/��n0�h��z] ��Vp�������uE�ج�=z"��u=�J��$o�1�U�m�RjP��t
lWWŲ+��Y0�A=��Jq��čR$t�7��~�Df�*˄
�q \T�be�r��o&�soBN1���0��Y�WA���������V��QD���;�
��<�CG���M��O�[���$�Ɩ�q�N��_{�l]6v����D!�b�]��Χ�ޒП6Pٞ1�_��ɚ�� ���������_����Kl�Ю��ǀ8��t�u�H��?���$��O{�� �ڎ!` �*�o���M�7�h�o�#��+�m�PtZ�as�̏�+�_F�S�pq�`�g�v�pߗ�l+�Ր*V7j��i'�4� ��L�	d����f6`V���>���Mp��#��D�N�3u�h��2���跼h�j��(������Ů�FO�����=o��|��0j�z�ۋ��:*�T�v#��zV�K��o'q��ӂ���y3��{������wt$� ��.��&�H�L��\o�����R$3�t䬔S�]C�I&��fOAn�?�Sb>�����"ǻ�'6F�O����@�z
3_M��� ��a=AӤx�a�5�d�����G_% ����գE^m�؏CF��h턧;F9�*J���b6N<?��K�=����/8��)_͸�ŋtr� )��Am	G��"^<Q��$�̚�	g��{�����i���������C�qk��1�_��1�1X����|y9&�[�)p����7�n�h�ƛ������0�����Sџ{�nl�-�S����:	�q�g��'����a�j��一�R1�Zn�WT���:~ri	�g��A\�.nw���H�!Z�w���g�4���32�&��io�.��$Q��TMsi�?e�
�����4mFgW����9[9R}�P��R@R��^5�����kn\)[Ҕ��5j��^+)i}�a�wo�����+�YA[û��y��x��O���M��Mp%�$����0�'��L�Ù�˂qR���͑� ���� �����)�yd���~��@ؒ.���U���i�D\t�٭��:)3J�enA����[�ē�e��߇�R.z,���D'���,c�#����3BBq�N��%@���\�@�`\��6V��3�~�=	�*�3f^�T�v
ah�>�v�O�Kވ�B=�Ȼh���x��.EC>�n�b�6��]�:B&�?���,>�TD<+�7����x�u@i�ʦ�k��N������
��	��}Jڸ4U.���/B�W�iD{��]��A~��,�gι���#�3����Pn�h�+c����E����/}�����*!{l���>G�@Ș]�,�.���4=k�M��rU���Q�ֵTBp�g��	�(��+�>���)���dWs�D� A��������NH�d#���.[DNy�B�G'I���:���~�E�Iq!n�Ȣޤ���"3b������4#��U��8�=����?���]UC6F�Ax4������(r��0iXC;�����g�g�W��77,@��'8A��Ïm;yd�W=&�'1}6����_S�F��i���5���
�?�F	����S�B8��w��O�C�9=��&�q��K�Q=,���*G%��T��{n$�0�e� �4bǎ��f�lf{�.!4세��fWT�i@s{�����jJz=���x�̵��y��V�P����C����ҫ�s�"��B&��y�ď#�\O���̛F-�W-�.�-RD��r98����ur���`�	���Y����~�SI|��N\vcI�-Gz�:�:z��+(���1�.���|�,#��f�!�	�pN����C �H% ;���+��������� �u���,]iO�����ih3cq�=wo	P�ȕ��=��"t��ԟ�A=BL������3d.��ɍ�`�Y"�������T� �-Ab&�R�]�m.QK���}�}������l>���X���{6��l�s]mr����'tg�f��=���y����#�%��W9�	#��HZ?9�䜣�6Q�6f���.+﫬��cӚc�v�w)`VX��0�N�ҿ�j���sx��_�`����8�a>+����#���(�������3�� )��j�t�K�g`�D1Y�hp<|T*�� zJ{e��5tm�xY�@�K�s��5Op�������.�b8)���M~���E[��e�Y�`y�yn���82e��UÀ��y�}��s�^�$���Ln�Yr�Vʻv\P�Oj�q�9�����J/A=l5�j�q���#r��F�g���S/��D�mn&η���z]���m��67VSb;S�_�l߽�&E`�'JF���]����cJ!����Z��	��5�^�3�W���]R�� JQ�亂|ڟ�Z��T=-��`S�g���XR�.�J�"愆\����@�����u�7�F��	�����(^�~�������؝A+%9�9�$�h�����>����d[�u- ��;�ٺ�v����	�:�.3]1��^&�Z��9GbK�H�A����Nn���yCXT׻�����Y������b*x,�0�S�ri��J.�Z0޾�X̥T�"_]Dy+Z7a#Vyh��̷x1i�w�k���*�WMO�ʿ<�� P,*�'*} �D:kBK�بQ#����)�-��g*�a�ك���^uk{��EU�)V�Ov��d����AƗ�3� �e��C[��E-�A�)ۍЂ�G	M��b��Y4�n�� ��k+ ���yN���5���%�T��Mӝ愇~�Oc����a4� ������%��g�CCN��:>���u>��ؘ��+���/	�Z(�����E����;�SA�3��kc�h�37�,^:���a[��7I(�q��p�ݐ���qZ�����������t{]��������}GV�Y{�e���t9 x�MU3�;Jn��z��_9�c�}�r:ǯ�y9m�_���)�h�_Aq!>�9&��50̭��>���ֈ�6�r�����:$~Bi+3�G7ö���}�;����d����������Sb]���QVI1���J{^���ʜk�\'�fp\���Y.�M�~��K*hox��]wY���*&�z�</:��X��zHk[���%/����X&�(7�\�!�}�_�x��Rf;,��FpFz�ϫceS`P���'e7�_���,�I�*�H2S������e��7*��9H�٬,���W�#3���#����"@��f.�0x���Y�x�񩥾���S��(|	��G!f�+���h�}����h�j�>&L���u]9j� �g�#��^�y�[J�B&��r p�}���b:M!HL��k�$7���c�Vť��S�dRc�����V�����^�ί���*�2=X?���S��kˬ�)�W��J�̩��2N
X�ʗ7U0��%�\!�S3�"[be{�=��-��NH^���L	óۻ�q���]y�9hO�UU��b=}������_k]��[p�ԛoşy�픐�`�2�Ρ�C��:�vnhyHŢ[��"�o���eK�WJ�;�}l�+�dQq� Ԣ�:��F���d8tW�R�
Ђ�º(��!�B`�R��W����Ëϑ!��Tɶ��Yo�K�*'��Ni�x�$��\e�d���Vݙ��8O�YΙv_�g�#���)p�R�Ѽ��)�L��%8��Tu��/@X�"���|ӹ�w�$	�=$"��й�ʖ&�%�ĉ�F��� �Xk����-i�
A{�9��?�j�bCn���@���[�|���5J�"��	�޲e�ݥ.�Wn���E�P1����j����ӯG�p����|��C�|�!k}�[4��O��md���"���J�5o��?�:: �$��V��Rg�_0K%�i�.�E<e��\����y7�D�}�۝	�A��g��Nџ<���P�э�Y��;%��z1��ธk6�hr��!��x��+a�N��i4Ѩ(�����:b/y�ak��eo�`)W"�dv�m����y�sI![c�4!��sq��̻>	8aZH�y��i\��U D+7۔���JQٔ
��'��^���*�8`2 ��rQ��s��M`	H�m��� ��bߨL�G��6�~��&l�4QD�EI(ʌ��m��]w{d�#�K ^ZDj���?�?�L��1vfJ���D�q����UvDDĜ�{1a4%��wR"*��yy=��U��#a��	�%��7Ζf��ŁFዼ�}�ai,��N��̦- 4�>4FK6� ���k9��6�]S)��!�˖m�_���M��FbDn�Hcu�,�0�<��[ ��1���"pYh}T��Ml���߇/1UF`?YH��qה�3Br��y,����,x�g��t5c���y\�yȏk�0��b��mU5� �R�
�U�C!�2�3[W	e�lLR����:`H���=<�epT�+� .@�3-�tv�$�ڂ�/���f�$ �ߋ��㗏�\�<9a�U� OUq����-Q�!X0��1I��0�w��n�$z�4�R;
�7ƍ6Sި}e䳋����:�y��	�cq� �ȩKH)K�/���>�bIt@�н᡼�j�@�Ý��F�����g����9�/�ղ!����~�a�HK �0m#����;�io@���\z�5���׊���[�g��.�
�����2�hF�6�yCo3�4���➲Cl��UՅAå�#2{5�/��N-mWK�\��S)#/D��^�m��APy�7�D����wxOg��Wг�V{���v�T"L^�&TF)�J���,Nz�H,�����M'��dX�^&	��U���xY�q,����\<9O���&��]���pC�A�M%����������&_0���D�=� .���:�h���3A�ſ�l��I�������j�8+L�V~�{2|���)� A7$g�%��R���m��\��N�Fv@&̑��vŴ1�ݔMJUB��EB�#.�۾�7x��F~�W�"� nCLu���k�l����a1�!a��[m��J"/��;�s~��٣��§JEy�3��n���[X�-�T��� ����i�-A׊�)�tur��`S��T"��IIg����C4?�EW���~#�gW˥�D��7$�k�m��桋�Y����aB�>�N��t�Y���r���Qx�U����͑�7��K��xV�t>�R�����(�!�H���%�Ԯ8����mp6����S��׶G�vI2�@�,��eeҺ������oĮ�.� �ſ���*�r��:�\uI��;j3L$M�f&Z�T���zB��O��Jt�?���Q�x�~fc��\�:�1)�WH��X
��n�8L��:��/B��F�x���K�d��^`��b͂d!NTe�fP��R�+:�e?6���sO�)�~D��5��Xg����pe=����
��ڄD�`�.�:�ƒ�㔥ab�s��Nr�P1��g9Z�"��6.�-M6��˟㣫��Y0���z
&w7��M?�إ;8�����I��s�@�矽���Z5:�u�)���M�g�J��K��
!r˾�Y�dDr1hQG�>#�?,3�ס.:�)�����-hAk�6�	7P�C@�*�|5`�����C��6A1y�q�w?� ��VcH=�ff�j)'�L�=��F\�HL�uw搏+}��|7qV��M{�Z�E#[8�ĠV�\�kx�ɘ�?	��)~�Sև ,q���dkNg8󆶿綇��f��;5v���1���-<��S�o'�Vd5��n�}������seEHYB��M��C0����+$[�U��	���Y�R \2��ca[�M+�)}{b�gxY3vA�AR1:�*���\<<�\hѼ�v�gz�&5���"�\c��th���+�?\��*ney̡'񫩽r�m�c@܉�I�ޕ�+�~�2aW�Ŵ�%��SS�%9f����
?6 w�,�x�����t�p��܅J�B�-'bҁnRs��Y���	�7N��)h�I���y͓���	��ʮ>	�	!wO�E��K�̀kw44�:T�����`9�j�:�W���P|�V�즒�{�W(Li4�U��#�������`��k�
���E�M��z��M���[|q��ƌH�ъ�iv�km�%�K�u,�Ok}�I����R�h��q1;F��7��J���eQ����xH�F�@u�8;8�WI���YB6�:�2f�[����)��oK�5�h�����P+��>�}Oؗ��H�]�9j����+��Y�i���.z�Eʹ��,�+�G?�Is)_f[ՠ�u�Qtz��9���j�ǡ���M�Ư��yX�;�����7��/Rc�������V���_��0ƯQޑ���c�fg�u�$�ʼz쪐�����f�g���b��JpV���xn{x�G�L�*�ˆm�[�!���0!n$�B䤼�:̄����"Ɵ������_|3B�=��a?~�G01g�.Z�1	�KTdN$ڋ!]�T
�����)1�X�;����<%�X�(HfX
�)C\O�c��榊��e5�^㦯��ՙ=
��ZO�B�i��Qh2oϗ�-�V��D�X�([�;�)��r�V��~���']����J�kˆx�U����R�(�5�w�K�ś��=d��`I�\B=��bl��T��9�Lo}�`������ _�A4������C������4��k�C�ԅ��9Q80�7�Hn�{��=X��*�n�l^�P�
Δ���/I�)����5�\�[4y�I�����/fĸU��d��7˧� ���[l/��ZEF��8���a�x���8�%YV�b�,��8(c'������E��14f�sU�!â
��ok��N^	�8fswo����n_��ц��X)���ag�v�;��z�8�o�� �ܗԉfٖ �D��Su&65����q��,��<��{?���l�FV�_c�/���0b��6'�N��޾������xwT��&�bc�+�+�? ���"Sb��X��TSɚHd�"�d���q�@���'86�¤��\ԕGk�r3�~�)
T4\|8�vi�^X5��怯%�NɈx� ��,?��ိR�a�N���J?{�sg럸JF��&���	s%�(�X}�ԛ�P�	�S2�%�UOB�K��}��U���F�	d��r�LJ7sOoN�݀������\���M�,�^i}�vH��x �V#~�Q�L4"�`�ѲƟ`Z��ୄ�Jۧ�R�~�ƌ|z��tB0�!���0V՚��OzlE�i��6K�`_�X ��(���=_`�T�
�	�Xۅ����]�]�D�IJ{���Jh,�J�u�G�J��s��o ��p�H�C+���:�B��z��Ld��6���t��r��θO���۫�@����+ʬ��(䩒%`Mf��z<��Fװ��2�yJ�� h G�E�r)����O�Ua�-s�qC@���u�5�9l��/3��<-��Е}ʩ����ӝhH�:��s%��.��Q΁�6�F:�g�כ����c����k����pפ���Yǂ�(R��F��ak�`CtW� �kz��b�z.w�y��hP�o$80�d�����ku|�"��*J��X����}��c�S���q�f`��[�#g��6��k	b�pc$*˛x$N�#@�T��*p\6�]�)#�v�ƀsH*NEi����{.(�{�GK��#^�֐1Xx�
S�t|�(��t=�q�a�K�c�)N��B'T��\:�v)����2&��N2$��`��+���>x�*�����]�[�'�¬��G�s����w�r�ޓ�A����D������r�~�I��N���P'�f���@ �/RfQ������6"l٫�_`'�kI���Mz���(?Le���jc���|ll
ط}V9��5މ�^�:�vZ���&��o��+��ƌmxqr��:E�qHЁ���qLf�(�_�mi���ߪ.���z���e`Ĵ���3H�b�O��̩���Υ����WS4~ jSi���'b!d��D.Ĥ`��	�����w��n���E��p�>�G߂�ȳ�qَ�޳���W���)��fNF�j�g�&+=�5^����q;���B#<���ICGЅRRMF1�\��9�@O�sϪޟ\��Oٶ�yA�,�GGb��Ɠ���lJ�#R���e�wT�c�H��������ع�>Hr��P���As�����'���sv�7���S$W���ټ�=hG��2������^}Ᏸ������m
�\��>t���T�'�8��>ū��s���������>��()
-��B��Y^TJ����k�_�hjup5��m����i�!%p�/�Ի����ܮ���J�����U�l$�xA�o����ۢ|K��=�'���޹M��w�_�.rdW�J�ϯ���$Cf���0�D=)�ؖ��l�'�~t@E"���G��D�+`���u�`&�	��m�gz�H�
B�:�G�[o���������H�m��d��#��3hU���R����^@��c	��EY��o(,����^�RL2��>;U��\��h����d@2��QQ=�����}��ϸ%��'[�Q[��%a�N�ԫ��c˞�3�$uc�v���*5K��W=N^�'��A]3ܟ�$1�+eYΚ�k���Ք� �f��u��z�k�7�Ne5�g�a�TW1Qq8��wCcm��ŧ����V�>��y�g�񛜦7oD��Vw	��%y1m��BKk�[���%4����V�������Q�V��s��B7��q���8|SO:@9/v�ĊÂ�TI=��56�*���$�I�tӓ�_�ڰ�e˙�����Z�M��g��q�,|�*#�W�"J�����%(`
1)����t�jz�83�d��M��rM����K H��2$/s��X��Bh�}����W�� Q0�_?%��ĹVbՆxt��lQ|�{)JI�bG����[=s�'��L��Sʊ�fT�BFk�j�w�%��hi�'-55����1j�o�?�X��4᫢�|}��;�cJ�I���aS�]z��} ]{�l�m|W��y"tw��a�vf2pk=bKpYtL�z&	�E����O�?�^�Ъ�L{\A����\T����x����j�v�c�Ν|�.��V�\��ۿ�Bk\_Y"���_;���y�q�qF�E������$���ג�a�U�L�O���<NN�N�-c%�K�?��r?@��!0,g�i���e�o��g���t����'�Ak�G.mP����y�p�hD������pFhW>�i6��ju��{Ζ�_�ʘ4˱\��Av���g��"]�#mG; V��n��	?cʃ|���K fN���<��3�3���m������*�}�h���1r��#�u&�U3�-�ߑE��Ǒ��O�{n����0��a 7/O��v=9?ո�|2,��'¹�%�>~�A֎�~��� f�}0�à$���#���C���U��n�҂�&��X,'fDҗ�Ҝ�'ƽp����%%Z�����#�V�|[�;����۱�nI��C�:�g����P�߰��A�|^<�K���~�`��ym��SU�{��^[�,��xr���:�:4ǵ~ށ֗8���.ͰFe�Dj�M��n��d��:����\��[�&0�K�#��'Cj<{�k�'������o[e��Ӂ�e��7��)o.r�b�3*��a�˻��q�7�IOmjބ�JU��Cۿ~w������`*�@��:���4��ę����z�g�Y�!�TA[�Ou��L���/��j��c�����4=��qc��3rĻWJ�,�.���c��x���u��GN�%�����	�C� �h��ȼcE��� e��Dsr