��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pgꍧ�i��;C�q�F���� �Z�`ڟ*]1�.��=�"�%�s�p1�IW��x�۽��_R�1�����L�ޛg�7Bz:�Ǵ�U�o�����A����cw��_Y<�%c{' �R2/E�D��ڧs8� �k�
��.���Q��������ϰS��}�&�f�"u���R�{`Y[T��>^U�X�G���hv��$4e�I;
d[�G�u�9|���H:l`�:i:i9��z�%��ϙ<ᱮL��l�<�6�jH���q����i�N����Cl_�Gޟ���'|x%+���J츈���[F����ϝ��@�����������]T�>�5h�O�-��6!�5�M-SZ� @�5%?V��*��Y��|1������|�f)�A~)��&��S�nTf��R@���b�F���n��F�0�&T�� �Ql1˟N��#l�{:�7�WW~C�J�aw�_Ek�o{�CE��(�fP��C�����O�i�|h����������/��ݚ�|K�[�2y�Ku:/c��D"�� [��'xa>[����wyl]���L��o`]"Ӧ�Ɓ�T���q����x�ID���Qm}\�-���*&1y���H�9���9�3y�{ �	�ǚ�4��a�ɤľ8�"o�k|���D[�T0��<��j>߲��#N!�,N}L����tOb��A�IDZ`A��QG����LuwD	�ez�C�|I�[�T�@�����K��lv�;����Ş����wfQ͉2⤞X�9E�B���7���B�c0��#��$"	Q�E�BW-��v���4�H���O�������'��V�s��_p|��p��~\�����9+|c�T(S���[Y"o/ї��Z�2�9~�-+�M���0�M��\�2�v�[ۉ?̾�'_xfx�7�u����XSG
���Zf��8K��I#^�����6�ӭ/	��h��f�P�ƻ�/�{�J�2z�����l��J������V TL�d�s>������Ki�C��&r(��0{�5�BPdxˡKvׂ�f���B��Ey��><a4�˻�Z]�L�4zõ̽�N�&��0�|@��h����	f�i2qe���K�1A
k�ɜ��N��,�� ��O9>�E�t7~`�ř���QEHt�
x���=B��F�{�3P���#���Ŝ
 {�r�{��@|����'+vhU~��Q�V1�`3�-q�x#��[���K�+C��X+5���E^�	h�� ��!�����au0Y��/�ro��ʜ��ؿ��]wKǫ�l1��œ?����f�GI���-B�ۢ�Rk*�-m1�N�2���d��_+���U>ּ�Y.8���4](��p�	|�9���;��݌�G.��`�w}�i�0�_��9/�S{ȫ�5��7t�@Zy�E��Р��F�����oKΦԢ���<$;)���l�Z��r���G,�;bW��Kct7YpBbA��VHIp���]E�?��nydĔ�G%��k�	�#\p��ۢ�����G�)� �<�`h������qsY��_k0r��(b��0�'�q�șݓ}��"�����Y9�lr6>��h�ty�`���Wu����6ʶ�f��i��:�3;��~��r9��f-T��#�T{���B'8J,&�v4���^�@���<�@�r�ǧ*E�mRJ��0���娅u�;?˞a�y$2���u��$��(���J��v^������~�_�P��)�.lr�v�0�x5g����.�e� � ��E���rs�������M��I���B�ɒx��5f�r�����e����M�#�o�1�V~/�l���i���:!�z\%U���ҭ2,��I�{�z��U��G\�?�d���	:��� ��V�+����u��6�)���V�2��������%9�:oL�*�[b1��hO��p�����}�+7X���ܺ��7��W&��?���Aeq#��ף������*M�]�!�m#����������2�*z��n�7"��X�����]j�l8:P.C ��A��f+�!^��zI�G�����W��D��7*'�>~����,�E^m���w?K���q�+efX�%^?���\�6�薨�����+'���By��\�S�Y�����i��x�����[�4=���X��1��Io��r�ÆhiDJ_D[�=�J��U��b	��H�[ ?�2���N`��e|��9*H�"�W�Q�k�x�5v��)I& �oCH�a.�<,����D�A�W�.�J̱�$������A��.`��]�z׬E��Ḁ���TGG̯)�i{S}�e���ǯW�ӆ"Q��g�⻨x�K?��R�vi��6�X5�6�߶�6X��,Sҧ�&��O�nE�tP�.C��e�<D写ϲD��eʲ,+� ���\^��ؾɷ!�g�e3��y ��3"|͏"u^�#���� \-�c�Y�v9čahm��!��^)����R�(C��,�����0���F�S�D�=�9�"�H6�^��̯���?g鵁�::�,}+t��D�@�+���	g�d�S��Ki�=R
#�j�����I(~�O��t�w��
ܸ��@�h�uG����{�"_#\ԙ��c��ypG�#�1ܒ��`.�^��إ�����N)!�/�g�4�V�⌎�1�P�Ե�W�v��҄����
s���NDe�ۄ���j��{��DZ%I�>\|�<Q>��X=�����ŏV&��	gu=D�Z���|�r�oԝ�HQ�#o{�N�j�_�47;��d����@K���B9G~��*
�9�a�Q1>�'�$n�/�
�/x�=�Ƃ������IH�s"���m��>σ�	��!Hf/��g�#eS���)�j��sow/��ч�kφO��	EA:d�~Fe�=�}7��1+/{~����N�)9����H��h�@�Ҷ��UE�J����H�?�#�l�R�>(�(hZ!@�<��@���N�s��2���@��[7L9+yCr�4�@�_���C ��ޑ�����l���OtG��D�}$�@�R��PV<l򿯈����-/
�^ъa�70��1/�p��W�
/�ȗ�� �8��J�f��L٪����^��J�~ %#ɫ�Ķ���C<�
+.�R\�+|���i|vLB�n27 ���C�jf�2r$�v�g�ez:J�vf�.����b��Q+k����䄉Ё@�
�8��.�O=����w��k����-��7�M��=��+��*�8���e8����ԅ8���	�i����PVBV���bA�s{���%�$�EV�;����^�_ǽW)Ú�
3��@���S�����m��$�npOt�R��D���g@���jW��O�+�� d�OJu$�TT��i�a��s@��x���p{�Г���8t�<
�E��^��=�"(FJ��Y�A����p�`��aT���մw�C��;>#��3���a�t�hl60� j2iQ2��g�̢{@�����32�����G�[��[�sk�F����$�x]���f��R����@�*���wS�
./�.��]�۱ϻ%�]�L��_�.z��K���#Tڿ%ā�\@�z�ߚ�T�HXkK��,��z��?�M���� �~גʐ� �ߚn�J`���j�x#���'�`�rP}~�=��0��&X����{��Vg�p(K���*a��v,�^.���S��`�wN��ݎ- �i�j)��J���K&�;����h
�_&ڱh:�'�g�����f&�󹁌S��o`t*jߩ�s^�٤��>&g?�o�iu<_��'ܢ;Q�^� ҷ����k��(P��@w��9���㹑a��/{p,�K+&�e92��V2}���RU�_��(G8A��.Un��/��踞ɏ]��tO(�xB	��\�q��n$I�W�����R��m�����eW~��!-��{�g�׍�_�Aq�W:p_���0`Z�˗�B���
��X�"���	҉7����1u�D�����ӛ|��p�����~n9� ᎎ�,��@�.���c�Rp+�/��݂�ZlF�0�f�.��*y�ǚ�ayX��:[	�É\��YbV����e1��AH�)�ݟ���_R�m��6�H�Ɋ}�R1"x�c�O�Um'w�����l"T^z��)���c�6P�����>���j���Zӄ>�A�eK����
ZV)$
Ć�X���t6�J��(��-R(�KW;8�\ݾ�����پ�]�@��N�'I9�s�,���鯷���������G���2�1E��HЎ���M)�Ы(m�Y�O
�j�Kx/V����^���5�wr�4d�6�ƚ��R7x�U#�����_����S��N�#�^�ym���t�G�[�h��*�`0#)�	�=�պ�R�+Id��B�	�0T�H��6ٯ��pFJSѡ�n��u@9��*�#w-�հ瀇S^0�r\�)�ehy�u�Q�Z)a��%_��r,�|�2��:��oO͡:BB�_4��Z�O�f�7�c���:� �Zpiǡ���0q���O���co���
�-��g��J�ȣ�<AEw]�&���ėӎ4 nk [��>~��.�b��T�E"��w��זb��� Ev7�xPAF����A@�;��'#@�I�����Hbb�����!�a�8AE��90��댧�o�x���W��n�6v&��Li�ho����b/���z���R�V���B�r��� g!�fm=�)�(�Q%��KG���?�zEO�cg�E�:��VxT��h��A@):��G��p� ����8 �3K�4 ju_ V��0��AkQ��L���r��pR�WwP&�ty�}?��Q��״���� �e>�x�5�>����o��as���HF�зL��!���E����^��(@#�X�!1�ҧt�26�^�5a�GX��{����n���<cc�Mw�R�g"��Wg�g9�f�jF!��Z�LB�Bz	k7��N\���Qu}x
�� =����(�]4�,šJ,%Bc�é�0T������\ʭ�=�\5Y�
GI;!z-0?�Q����ഄ��An�΍� �(�L���?�'���� ��(W�b����^,�3�Fs�m(#~�ݐf�4�*C��WY$��ެ�D�a	ac�s�_N�-$�H���-t,I8o�cQqӵ��>�Y`r�2������3u=Ƞ��^f�ڀ?��dd��o�M]2�H%�8��X����j5��޽P�m��Ft�ē����� l>w)��?3���=,��-��/@���J��
���u�:����O��^�G�e�]HM�)a�>�Te�4� P�������l��ZUk�(�C�ypS2EB���V]� j��Aș��7���"תݺ�95 �|�U�_z�kג��`b�X��X����/N�LV��5���Yɳ2�Ľ׶�<�Q���*�PW�ζ=�{O�f�����%�x5A�����mj�`k��A�3亮��tN�3e+�ט	�L+m���ֹ�4���<��b� f���M���y[���b�km'��t�_d�dSp�G*��������v`"�F��}���@r�����[�b�9zB�*���kF��l�q�����O�@Z�����N$�jm�Ѥ�,�2
|V�1��t���W��3j�+��9x�F����-������N�_�2�H#.Q�������ʆ��p8��p�l��܍[���Z�[±�L�!fM$GB��R�h&�������O�bi�,����Ծ�1��TD������+����UU�)��_8�Up�#� �/��:6�*��}4����Le�&-}"�#t.�K�E�������e��Z��6y�{�r�z�[yV@���l������F��C�w���a�ЫI=0�g��?��-�#R��`@�������,�o�זH$� �D2��zBT"�g�S��v�%����Y�d|��!S|�pr��R@**��S։�q�\*l��_e���~�ϴCn��cf�P��W�e�k�=�����s�g�ږ�ke�H\]�L���ݓ����,�`J�|(p.��������Z�G�C-�.)vT�:r��Z����
;tTw
�W�fYz�NI����5���LC��3 V�S�`O�MM�E:@���#��G���:
�^9���U��!e�h`Uת؃y��(?��+-� p׌�=��vR/���"-Ŗm�p�.�'�4��J�V^��6b�)0u��j`�(�
�ۊ>�ae��_O;h�٫�k��6��T�����~����2�{+���2
��zn��*)+�_��@�Da�C��G����}Ei�ۿdmۢ���nH�x2%yK�͜��I�{nf��$x!���y�&Y�����.$ôb+h�1K���U��
s�,�/�!�t������| �'��\����٨z��6���	W�nh��v�0ٴ�ؽʬ	nb*���{�u0�~�������mf�E,��K�q�����1�9k�w�C�uI����Gr�?a[��4w@��£���m�>*u���Ʀ+��$ԭu)��5�S���V�Z�_3���G�'��X���!�7akj�W�E~�+b��d�;y��1�HI	p�{R�;�]i��%�e
�#P�j�G1[x& �������TS��-Q���D�dCD��Fd�o�������)�܋�0N�<5s$��kf`��w����Ԡϒ�tAI�c
FB��h�����2����K�v�d���*�@�}20S���=��ͻK!�أ�`�He�׏ )��]6����3��`5�X�KZ�K�V����o�3 ����u𣃷�M��%�!���� �~am���������lya��Lճ`-)bx ;�8�ߙ�,���9W�x����u/绥D۴%���;L�U!Ȫ�*���@��)��c*�Kd��r��1(���F��"�QU�U��3X|���K�$�+�:��c8�_|���6F������~��K����@3���,	gb������I��\z��)v����Klgƥ�����+7x�� ��uZ\N�w��a\��Q.�2J���oyE�]b�-��V��Ll�ZO���b�f�*h�^x����/FzP���۪�'Qso�FYM�5�S�4f⅋�J��[j�iZ
�@w?>"'��u���Ъ�̀�䬜�8�ɼ�4�l���}wt����>	��LZ���F�J��w��G�I �e��%(Iz6P�^�h:％�"/|q��߂x4� f�T�a��t t�u�3�u��Pc��?|���.J���亡��%UO9-�� ��Ȱ휲���5(/r�P�me���2�U���{�l,>9_dk:�Ӝ:����t�^��������ʳ'6i�����%-JÊ�W�䷷ӓ�{��M����&�NjZ����h4��7��FF��.jC���8 ���n���@D!2�yG����a�23SW�U38�MŴr֟�ʳǷ4I�F ���`�/���^��F=���q�D�7�eu��F<s�{�S�Q�f��&B�ç藌�ZH�
X'z�Dَ�5
?a��ݥNՉl���U�r���e�N^'�v��BXQ\ҩs��b#���&
Ҳ	�#O�Ģ��](O��'�"��i]]�@�Gc��F$��D�"�l����@�r�����a�^yY���O;`�˾u��y�P��J
��O�����No�3� @���αm���ȗ>`�!|�CK(0�<8�;�g�/c�< �Et�<���دXGì��(4��R(��!?�k�sA7�v��Z�R�عѳ�])᎝P|���-&�9{�ʀi���O
Wկ6$1�hQ@���#�Vޔ 9�w����平���]�hLx�.{�2r��7~�Lp��ҷ*P�F�/qD�e��*H1��]����\ܒ�}��w�5nO���}ʑ�!ʰ=������q*�Q��_��J �� �hZ���tK7ނ�ošV9��y�M���:����Ȉ���XeD��&�m �{�E/�����'K��65�'���?�${���b_ǝ��������?��k@���%�a�Z��C�%��$�dXO��	���t�:+�!4'x<"�S�,y���8���o�F�PђJ�W�בe���w����9�g&�D�⻐y�~�طE��v$M�fW�o��W�o���ǯ)��;��v�S������!���_t=�&L�⋴��&��˾������ Ϊ����d����<4�Mj'��!{`%�����t��Su��*�}���+��}�p�$(�Yo�G� ��57��L�4_Ҥ�	P�q����4Z[�W(w䎥v���ťխK��	n+Fi7u����K�ua��&��T��1n���S�:S3����JR)]3v{5���ҩ,���
q���t~�U:�3�	V'*_d$���-�ӿuD������,.i���q�!��7��{�w�"�1�[����jv1�>�E�2J�z�oǗZRp�B5?�k�Ȣ��h��������pYkp�m����s]l��`���S/� [�=;�/y����9�:GA���� |�Is2�*[�{o�p~�C�����t{�]2N����_8VHq�rX�ŏ�����7��� �?^յɥ|�:E=���g�DHYZ�Z�/GnD�����y�X���KP��t��#���t) z]�4!��70��˕���ꟸ[Q4�_���)`R���Y?�y�BSR�')Zv��'��� 1)_��P�cЃ.�^�ɉm>�h]��aKS��*o*@K���6�:ߜ��E��F��?���'"n
 >y�N�z�CQ�cK��p�y�&��ˆ�$r��@��m�Px�8�h�������Z=ECBE�dGs?�Ԋ�.��-���D����52(,G>���F�9��)֥ꁆ������X���OqD�>b���;d��!#}�$�a�lT�C*��sz�$�l���]�u=��	���Ç���\���S-K��y�;�o׬Be�uz�� �<�"�Cڕ��sG�Y�n?���- �4n��6�j5^o!o݋�g��l�����c�"1�D6���[S����)�E1���"�̈́'�jY�G"��- :���i�u�XZ
y�d.�m5cڀ�MIU����W3� .�'����T����1A�M�ZeL��b�%]蔪��J��LF�,=3�6Do��|\�*s����Ӧ;:�v(wf�Hn�_��p��u���0ԑF�w&(;<���L�Pl��w�2���ʏ���[*��pE�;샲�DՍ�~��|����K.4�0#���z=�D�g�f���h�d���I3#?�v���>b����u������f~�LglNN��N5��zJ����h�����J���ȓf�
a	����ļ)uӅ&7:�6|9��Q��[�NF�������&�~�_q$V\���G�+:G��]Oe��2'A9�R�!��M������Z�#���M�yt��MDn�izb���w����b1�	�y��|@5+Q�?2'hU.8DW������W&��Z�	��S��	����9�˯�������m[��"Q���(J+ʁ���<R/��kj�Y	�~��ܒj�y��}����p�(1��k38!pr�
�<��P��9gK'��g���\t��8 )P��}~-$��W�!�X$�Sv7�mQyb�S�3,b�r��>�cي}��Z<k��g,��?8��A�f����pF��8	I1;Ux���V���k��uq��U'%t[�S?��~&a�q��G����8��z��w���ar�S�Jz�L�ua(}d����������Q�Z���	2��=q�_�,aé�=~��u�1GC��7��5��#�Uk���C�8�58M�� ޲�?��}�2�A�;lC����`��X, ��<M@\ɤ����@Jς����7��;��1�	d�O;�L0�q�����&v5��6��b�" �Pl��������]�SA|j#��������Eנ5���#���C�U�N�����yę���s������鈷D�Ω�#��`�]o��A��$�U�F�!��P��Z��,Aw�$�f�n�BJ D�utR (�㳣]�e���ER����Y�J��y_E� A����<���s�%�=������h�>$�4�����k����D0-U< w��J�ܝ�g^S�W~�,�W��F�H]��?��[
`h7��������[��Üߜ<����L���<K��+�b~S�+����_�t�E�o>]�6�4��JdaGV+�D��S��)��e���?&�}ϭ* �>�1���!��C�tnK�ө�!�xV��{~�7����8�Ջw���ROb�E�S�j:8kk�3�|�
�x�
����YLU��4U�T�|���%Zw�-�0��ŀ�7�fWj��&�O�)�7�5��+;[�����:�	ffZ�M5�ǂ?��e��)��T���c�s3$�$�W��j�����qV�X�X,�hl�I)��	��W�(��	Peu����`��X�oYI�].�?�Y�k�����nД����X�c�}�k��q�IC����$@� `Iϝ�v��B4N��6���rmrQp�%�\͊�3����\��@�ņ��LnN�hCݟ&"_-�g��W��W-�0���n�(|��|-�������"B��|��g&�5�F�`Rs_cK_�:�,U�{�B��`�,�"�A�� C��D��G�dJ��r�7 ���s�0�	E`o�g�����ϛ��CZP�`)�������ѐK�?%#���$14	]���4�O�vA�~��0 ,�}�-ט�?Ё���I�hH	���N�UT�PY	&���8�V��gq%2�¼��(/yOZYJ��,p,�%��1!!�S��e���cq}"�`�Lx�k���G��^��<������� ���>���^f����BjW �xIc.��y�EL���q"�|	`dاbӯ�qL׼N/y�C�J�Ъi�H�������Vi}7.J�����kRa�e��.E�_xE��mi2�B��������@��w��+;���j���/i��u���uQ~3�g�4�'㋇�%�'-@�A��%�S�iYKg��%�T9�A��q=ww�:i)��}�<�&�WJ���b����L1�;Ї^�G�*�����{�ŷ�k�U�c��q���A�Ʌ�q��Zc7�SW!��)����=����r���Wr&�{$��iyύ�ɺ-iΧ@9*u�.ۨO��?�h�,�tD�rȬL���,w�x��U��@�A��ZN�����+�ज�>���
��F'x:�}����O_�Ȝ݊?���d�l+����i��T�H�B�%�0����3�r�]
ʸAD�,�Z)�X䌏���X�Z��Y1>"Q|��ȟ���u�fW�>]Tl���f��p��_�)�M�_8�˃�Δ��!�B�Q���ܜ�v��/2��h�ޯ���슡1R�f�u(�^~���(^�ŔU=��;q��2a�;��ņ:����-c�	l'd#��Y	��#Ǝ�	�v�-�D9�H�K\8��3a���
�A6ɩQ��w���� � �����hF�?�fِ2��$�Ɉ��ẤG\����1z𘳚��1H���֥��{��}%c2�1y��0���c^�NSH�&v1��Z!���(uL�R�|����T���<;~��A�Y��a3wml1O;Χ�`Aa���">�o�)�����+ ;j������ω.>�}��SU�ł�а=_�bҥ�C��3��G�AS�KQ���v�>X�o�v��d��!c�D�U-hQ��1u��b�<�<{���hF�r0#X�W����R�o��6 .�$0�x[u&�)���o1�g�j�
�@���a��B��Ԫ��iIP17�1O}U��
�k�������r����-�����Z� i�v�i
 �d�xV6��8�����r"8}��� Eկ=�l�D��Lk$&�h�ssk~١���� ސc�>�Y4ʁOc1��y��O�8(��%��q �G^2Ϫ��jmUD�\:<�^��)��U5YT����q7���{�zN̄	[�.��*�%6�*��<���Y,�N.���� cQ<����g����	;>��P5��'���z۬��/f����� ��Y)�� ��b�Ԃ{{,�~@�����\��.6��� d���j��?�%s�_������ۧ��0PN$��w�YϞۀt�CQǙ�w�ԍ3bJa�Qd�5#rү�ry��=�(Yi�u���٢�WS�Y�S[+o��l5W�2����aM�[HK�t��i���T�;�d��㫦cN4%-3��
���`�y�)�j�D�,��v�Z��d�^�V'\/q]����M\�����O��x>xq��w�>���kj�$��.��]��[�9ؐ����`��6ғ��[rߤ�.'������$:��<o����J�������C���U�ٗ����d�`���_Zl�0J5.jYUQ�'$	��O��X�)� ��s��E ��S(��U9�7�tQ~�Xt���BT�y(�\k��[Yz�����/YQ\;�աT�
Pi��x]�����e �� P�%?��X��x	5����/=*�����6&,I����n=z��zbN����켨0[=�z\�����ևF;�Þ��D �]VT���	����X���F��v-����k���N�Ul��gW�ⳤ��Vy�Jdvg�?����"|'#+h�<5��v����-���1�@�/@��M)00��1C~��^�'��C���q����F\y��sC�ߞ2���Bۼa q�6���Z\��w��v�9	?;�AxZ��Ү��7?���B�@P�a��G�5"8��K���Vz>$�o(���o�Uf�\��[�E��/���a��&	|��b��[!_��T����w�}!���Bg��Z]`���YgQ�V� ���:�ƸfSd뺳
��<�*T׃-���EY�JM�к}⁧I.��ǆ�ֲqU��:k� s�|�@�"!ݐe�K��&9;L�vҰ�I�vBl�D{x��1�K]�w��,dx��x�oA��p���3�y@;&�Y&�Q8v<�@M,F�-i�Eq	���F��8���qi��h�o��<<�F��O����X��V�A6�=�06�Z�-Ƹ�8���)�r2�]\�DiX-���J#AFִ���[�l8�`�u�ϼ�Uu]2%tb\I}��j.�xv�F��Ht����ajzt�!�I�n��&�c��$ˢ0��SWU��b�ʉlH�=���� ��'��$m��u�Ӯt� �{8+�ȩU�$�/z��z�b_5�v�m���9�_|J���n��Z�>���6��c��hG�~�����C��Hh!^���Uo�����9dg()ˌуj�@�����Z~}�gtj�;�����.1*���@O�V��m �E�R���.}�4CH(~� 8���> D8&��������!�|�Ϣ~�/��L\�k�j��i�3�C��w�=m����~�S��;���
�����<4�Ђ�}�Ͽ�G��D�Bϗw}�y�6�dPϝ!���|�p3����[��91�!�WJե�ujڼ,o���a� *���gBD�Ǟ���]�,�b5�	�t�����+�3J�(�Xޑ9�m���?������W���r��n���T$8���Tq�b���8/��,I�����썠5Ja!e�p��E�h31�;	�M�$�cj�c�b^7�l����<�I�
��ڈZ?�s�u~_z> �b)F��γ�b��?{�w'Zd�c���|�R�LΡ�T�gĭ֒sD+��&L� ^��u9�>c�Z�7�C����ik������T�hF���O�>�� �8j�����}УS�7�9a*�)�8����֥�R�;Kq���삜;�=�-b���Ĺ���5B��*n&㧟^9�/�b;2ܐ
S��dС!kcںd5Z|��$t� {��9�\*�3�|��}%qv�{FU�P�s��
e�O(T��Ue�۫h�.�Nr���k)m����4Vk�Bh���?�<"j�zhtj$�����H	�;��;�̢^e!A���dt��{HŘ��|MB
� ⿗� R옪\U�Q�1V+;f���*?�?���L@����X�f��o#� �j�T� 
���)Ž��ñ|���`N!Y`�"�SɔO�� �ӵ���/��9��6I$W���.c�Y�v/��=�6����D���1��\�b�+)m�Ҫa�k�����Ο�Z�����O�1+u��=`�߫�"�6fG�@��Q���`��5C�^5)��z��� � �d��7&e��v{�G�Va{fu�GhTaᨃ2�,`?LB��� t���v��� �4_��F}�r�0������6��GB%�_|ͷ@�Ѕ&�QR�f�#^e&4����RSd����A��ʄ�b��٫�]���G˦}���?�W����Рj�`�f�I���@q�����DtҦd��΄Ն���Q� �?��֕����"�#q�+GW�6��:$!/��\
�X�m~�z��G�$�D�������ŕ[;Y���+l)a�7��m�y,I��t�4~s���-�5`�Z�/���&�n�����B��L�A& L<�n&c��>̡F
�Lc�7Ѯ�4m;�W��n�$��i�(s�z��U�<���,�*w8٬�t�鵗�ё��?Q1�n;q��#l�kU'��L���89ڦ�	�eY�54�4��N4��c���Z��r���y��T��-MwKL�Z m���N&f�e}�5D8,�o�6Y� ��)CJ�Ґ%�hH�j��T;*���<V	�8$��H-�g������$ɖ$�`�W��"��D��1ڢ�WΩ6��*uFr���ulj�F��/K������[��k8�4-]3�Z�6gI:����]�|e����sP
�����)V�Ֆ�뷵�9I����&��ڨbcG��2�B=y���� ��fE�ϑ_�ބD* C�I�.?��:&�k!�%5�w=�5n������ߍ�X��e-��#�g��M��e���H����`�[�r�Rw�#���J�=���S�Z�N�p�P���nX�ǋ1۩R�2�*d�����:� �t,�4�O�5i�z����ǜS�{�d�˅�Ekc���yqKiCe�y�����r�(\����m�&U�eT��"4��Z����63�����5e�A<$OL������95Kl%R�y�(ϥ�H5�mϽ6,?��ޡk6a}�T��6<��aDJF9E�ŝ�n��U��I0>�}�c�X�[$slH�6���E�h�|�=�����3`�Ah��D��$����b�ƽ���;�
q�V�!Ou�k��~8��M�q�d±�O����&��r��ߖ罏ά���2#>�{�#�Ж���_�3s�� �Ճ�ƫM�2o=j��ӗ{��K