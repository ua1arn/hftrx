��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^�u��]]��c���Nd�e�@Ѱ��iw6���=uC�Q�׾���VL�����EQ<gS�Jdq���<��;^�<[0HFI�W�W05��p*x��$���[��l]/�a�a�U���k�bS���c���;d�#�{7H�2ŋ��J�3��Gqn(Q�¡l��uw��:GV|����J�'[MU��0qZ!��*T�P6٫g"���(�4s�4�f���_���3���=�3|�7�(�n¶Ē��P��ٺRd�Pa��vH�r];4�\w����F�XX��Q�AF%\�#�eM�5�K�5˧־}�G�s���P����a�[�gƉ��銴6	I���&|*�g�(���`|�G�d�q�jz��2��I1 ����׼ܲ�5FZc��V��\�ee�!�"�ĉ."�,�� 5�ݕ�?C�P��{З�wPt*��@ܯ����g�/����u��N��1P!�F��R��U��\|z���;5���d���Ȓ�w�}B��5�z�M�����+S�!�
��$�36%�f��Q�\�b�Jr;�Gn��Ng��6,י�����>9�x.r��u�3vڠ��M���/�f�s`�g����J�9$��6UGV!�ʟ�7�3L긚	*�����i�5T�rY�I���G�ϐ\�[���ᄯ81��vN�	�I�\	��W吟C�!�OQǳ��Ҹ�?��_���蚡�違h��v�|�v�E��n��=�������ڏ��ma.��<݂_�����y\b�V��p�f���E���>8� �t+�x"�ݷ/�]��6?�>"I�R���u�0�����%kĵ���`¤	������e���M�aXy�z����HbG�	������,B��M�G��]�d�X}��H�l��n sPt>����^t�����'^&�.�`XQ�)]�qX8O����O;��EN�����O�"�GCu�XLQ+`Bow�;f5�m �?#n��.EV^���#�>?�C�����̼�}���j~�����KC��W��S��8m��m��V��_�L�o��@Q�wq4ٛ5A4�Y[��YWm���#��������~��4%�v�6ܵ�}!>��(:�F>��ډ[��jLVN������$��n?m���A79���~�@���4s�HD�@߯�����`b�UU˭dj��l5��yECY��G��S�Ѫ_I�8�����Tn��}b��r+��#��E�S�G�s�Nt�1�p7�v%b��ݾ�;A�rŻ@��Yj�-%B���P�Þ\m�������9�wdTHo�)�	� ������&_3�oN��9j��Q|����#1� < _yc�U�x9ZFB>��\���}�q�`y�69iC*Pܩ�(X>q�s��O����Ln���9|��z9��:�u A�+� ~ȅ1��uy^4YHۋ�����4廥�J�?����x������j0x��]@�$��"������:g��t��:9\/���Pn�^$ aQ=xZrj;׼�1pi�Ǝ=Zb� ��JKq�̦�D��^Z�x��V��)��{<�H�Qa��L@���v�浽��o��Mf9U�||�9h
�?D���P����-S��)j*�v'iiP���ej��8�GX�y��ig%I횑�1�m�&��Jfue�a{ڞ-.f��ɇ��OY�WP�g�	�5Ёo��YM�e�Y�����%A 1d��c�#{�g:*} ��7�I\*�����P2R�e��7��*p��أ~�'��w���9��j�^X����Y�#CϿ<z�m�s�ǿ�����'��v��#r1��~�����e�o8����-<�~Z��Аj<F͠%F��]���n��*��;�ByC���9Ȋ��j�c`@
�OR͟�������J��љ]��[�+3�֚cϬ�ǜ?[�+%�rd�ԡ��N��zf�� �ܮ��
i���r���Z�=��w�?="I���tdQ�E�p�\����+;�%��ū��h�:F{z676��ro��/s��޲A|J� �l�h�.�S�c� ׉�����zSi���'�TJP��<�ɯ��ݏ��ƚ��	=���m������@u��Nb�c�NA9yS�������٬%*�5|f>5̣�$P�#�I۟��dB��+w"�FB���ž(�+�}�6�^����[Ȩ�*B�ਫ਼_d$T��iR\fx��EU�}.ݷJX��ۢ�v�,�ݭ�J����Z��% �̸�}���a�'j�
����?��ۿT9�������-$8���]k���.:�3�b�5�/u�N����ݚ+or�W��L�V2��W�j�!�}�a�w�c>W��L�p�sJ����M�A%�t����ՓN�*�F��4�H �b��t f���s��[����p��=�!��KP)����Ib�!D����`� ���!��h���P��D�4�r�L.�$a�@zj�F�q��ݢN�(�xJ�s/1�DX����eM�>���&�AϷe���;m�M���1*��H�-n9�`���6���y�1��;�\������^(X.�a��`��3���k��[�_���BA!��ٙ�W����_�����mUUb���ѯ�ɬ[ +AAP�S��e���,��O��XR�U5`^�I����*���
]�V�xt�K#�J� u�����X��l
M��y���{ 5sPt���J�)S��|C�-�N�x�Б;Z�鄈�x��kD���5b���9����{VT�tkp��Dh�ƇEXҬ�L(��5����uV�s���󰐢G��Js�ęJ��SCR�h�<zp��pen԰��Xu��n>�;�A��A�Π�NJ���/���j(m�'��
�z�<j$z-Ɉ�WO��~D,�J��q������|@����b����Ö��M��n�����)������81i1.�~K�+
#��LM�z�h��X0Q�&jf�|�H�'�2����K���>���Rʰm�q��X���j8W�������*`cngM9�tѭ^z}+��_G�E��SJ�����NN��ף��~��s���w�rꨩ���WL�1�UCu�{�d}2�Pfv��ñ꥽R×�Yn��r2�KAY'��~i��˫�0�h��F�Gf�PyH�Nʻȕ����]@�[�6yI>���t&�?�\	�c'Uq������5S�X��
}�j@�.^�����,��ў���0��>��q����x����A��8��>i�U�+��1�K�-B�n념�<�Խ����ܠy'����>쪚�����d'S�M!�
V�%�<Ç���m�� ίjN 9����Ԋ�o��כ�0XL��:��e��Q1�=�4��A.�ѬY��ݧLZB׉�i�#4�����ꔎ�-�@��R�����n�u=9�lrPu�����S�j�.�ɲ�(se�s�����|����{W���U<��Ȯ~*V�p� ��9�1=�E�/�Z����!��w�Ҍ�>GI$+(�
��QH�kz~t���q,B7�Ec�6�q��Z��Aӓ���O�~t�S!��c�VS�`�𞐕��� ���/*ޙ�{�/�mnl����jK��%X�9�/Z[E���83�F�t�t�T}Դ���\=�C����]+'�z������u9�)�V_`�8>�\sn%Ģ�h�7 moV+��W�/$[�A0�j�s�$�vĉ�2pź�	=���~Z@-\�~b+LF�!وs�q���'��#8�B�L�5�2��T.AҜ3��I�1�g-$f�)Q�!S�y��ذt�mj+"����-�J��X1�� �5��^1�����,�����֡8��g)�z��m�T��M�<���{�M���I�黚>^I�t�����#.�������Qg�R�i2����E"=�Q��nu���w�g�w{�'���[Y�`��	d�ʃW��#Q߇�gKeew�߅L�=B�����ɦ�L[[��s!q�	-y���=�q���<�=R��|WY� "�mM��~`�ۇfu赣E�*f�+������E<���@�(�j��8���N��!�� ���[پ���aRJ�F��Xe	��U��L��v�I-(S{�C������C-,'�%�v��@����Q��4��]������Y'vi�4��U�������X�S2;ιL�>h
��V�31�ﳛ���;����8����߸=�ݻ��.�㩾��+���fC��";��5��J�B�&�=��Y�3{M�~Z�b�и��8�N�Tw���8.#"9� *ǎ�m��P֋:�8�k5gǟ̀%k�'��et:��1}Х��E�љ�b>���D��o�Cj�
e`rf���\�e��Kw���'��qx�өT���ք}��	�m[���԰E�N�j_�:���N#�/�r�ڀ���wC�y~��� HS(4�PɁ�3��'7�Q5m�rwG>үZG;6Y܃3ƛ"��X[��u2mћ������3�L�[���P> �bA�����DŇʫ�YWE�@^S���D����n	�D��?:�\"�Ϥw�N��4U����`͖�|���@]1�7t���t'K��Q�WUY˨@�����q���Z�@$�}y�������m$J�+� Y'J��x0	T�u���0���Q1>�� �v�?��-G�Tߍ��|ϯ�����<D�|���4e����s�@��]YRjV��"Nh��,{����eTה��$��|lu��O0����c�q�:�&�dЃ��+����~�ٖ���@xi��~]����#;k�~�^r�$�T@�e,�=�ul�҄;Xi�5�nL?��2�ˏ��#`�a��3"����O�"��?���K[�n�M�1ⱋE�:O*=92:���@Z:�Xґ,vdMަ���!�O�jt�f�9��+�bt!���2`E�'q�:���c(|ɼ�n��g��Z��������AizY��ﴑ�k1�F�zWS)�S8��u���@���Z�jʡ���G��B�<��e�"�Ah|sz�P~��o7��t�'8���n덆FO��B�/:�,���q�e�8CCP���}IC�t q��|���&v�Ȓ�]$\��Osa˚G�{�mI3���.|w!��E<#g~�4���@��i� ���?n}��$��4F�rQl&TJL��Q�y�� 7�ut�ΰ��4A�B��ygS�-ҟ1�ʭT���;�\]�����	�)���N����V�p�3�9�����1�m5� �|pVJE�̀��p����93h|7u{PfY�M���EE.���{����	�C���핅J��;�[K�����3���:2E�똄n16�#��f�D��	Ld�[j
Y�զH�z+�נ~2j��6%�p�e�y?2�굠?z�
��QF�ڙ�>sR����I���)��:Z�c�F�ރ%�Л�,�GJ��#�\p��Ȼ�&�ud���Ǡk���P4L.k�C%��mvG�5�Y�[�n}h�(�0�32ʕ�R7ɹ�j��h�iV�s��d��W�����
�>���4�2�9¾�zA�3��s�9z��1ޓ.�i���a�����L)����w�du�az�Ļ<��p�L�?��zj��9�"8�
hKP�+GT��9��q�xg5v���x=�Ad�[0�uW�w���VD�&Py(�P��H��.��}��c��z_r�-����Tݎ������<�<S>4�R<i ���(�z71���Wf"$��QY����������bI��i�(Y��l+��`d��^�ѡ;޳�74��K��m�<4�Ho�5(��{��?����ܰ���_+2Yǝ���E9~{��뢆}������ŧ��lD/q�$�)��>��0�DޡG�׷�&�$�3f:a��"�c�R�D���ǁg�P�v,J���>)1���gD.�R��1�rnb�S��D�ױ��l�櫈0�s�|f�w�9���ĉ��̣�kB�SՀi�~w�fi��B�h��5>��|h����ؽ�T���D�5������3�a;�6D�[H���B|a��U�ʗ���\(�ף�_m�|�A����8r�Tj�P�`|�#��j���+s��[8��{�8�%c��H6��ܾS��������<}���&�)�R����Y��(����.Y�\���b"�ZX��ڐkoa�����؏��_�����!���:�.U�����H�V�����~b��ͬ�OB���@�t�D
�m�vF�4΄[�v��@�(W�o@U:�H�Тx=��[����d��jɒb6�f-��k��jI;����o��A����xޜ�^�R�N/u]	�{E�N�����u"�d C�Ş��Ȉ�Z]����
6�Вl��.�i%M�iw�|�~�,i.��XQ"�4*���-��NwR_�>v錛�YA�*���Å��'�"�\�?h�&�#?Ͻ���J!8��p0��+�z���Ͱ�;�T�����`�e��C.Ձ+m��y#�2�5��}g}�_J�ɇ{�m!Ce*���k��i�:������9	��@q3��Y<l2�V���<�"�M��J7��Z	po�2ťІ ]�yc?�SEzs����X���������<�hG򅮇�������x��ذ�e'B�c*Pj���+�HE���Zn��g���J� ,�^/	k��aTk�r�~Բ���ox�K�Q����ct
ʈni|suM��7`����_D�����xc~�a�}Y���'�iX�.ʮ&k���3oҩ��P�4p����	/V���E�U�ne���@8-��<7���16��J�j?:�����K;JO#J,���0S_�Ȇ�
�@�������4�<IpTe�}׆�I�!��ѽ�\<=��d�2���Y�@�!��L��Q�y�{7�x"Q��(�5z�7���ˡ������!�"��q~�f�Q��l�<�E���SUp��f���۟�#V�q�կ�x�@!�=:gj\�)
�P�\������;�If��D�^�n�b��@��q�b����	�R���W���Pȗ�����h`������R8$���M�cj�1ʅ�Z�[��#P�2����^�/{�nX!e�\������0%}	�L�`�d7�K)'j����	�NkuN��@�
��l�b�1������x\�[1%tz��ؘ[�as_�7ьnY�(ҿ����]b33�j8�r����yT	��ّ�9(��^C����aw�F]=ml~�04���0�Z˥h��3?;�&Juj����,����VSlQ�`����Vjv�'���Q<�����Tb�Y;�ݽ�x&��ߛ|������H~
�>B�3;ʐ��6�s��qP�ݔVm<�Z����졦��8��
������7������wsv1�<��"�DM�<T���ַ���^E���7����9b7��Q*�I�"� �T"�A�:� ��^Sl*oP".�r^�\�ܚ%兊�3����1�~b�����՟U+�s�5.\Q�������tH�ʹu�x��n�|w�Z�I�h]��J�q)y%F-�'+qd�<�b�҃��T��'�����������	�+������M�!�&H�h��+�����;4~��9�D����
fB��c��6��݃�Bw�d� ���B�6S�-�W��ފID�E��]��N�1�w�n"	�&M�W���3*�fX����s�x֭� �܀"��0����qF� ?S������~c��n�"*	��x�nyN�
hr�(5Vnr�I�o⹡ �����M%q<`��#�$������I&uW�J��}�ޤ��H�~M��B�Q씣�m~g�Ǝ��y�a� 7�)�����S���v�b�M�e�*���~_�C0y��ӯ��b��� ��S|�	j�֕���l�Dj._D�f��H凘�T�����I���O7[�[�����-G� ��Fr��H֖}��Bg`� ��*ߣ�q`E��5k�7�1h����R�ǎ<t��u��Za�s����{���,0o�!�r�W),����+lߛ�I�ߓ��Q�-�8�Q�I\�I�n�B�gcT��d���7h?�b*��57lw�CM��x`M2��{u9W��D�[�W���������Ʋ���6����1��vtH?��]�(T�f4ŀF"F���sV�kB�!Z��8�a�S(WtÇ*B�ͺM�4�$q�$\�m2�Zy�'�����H��F��1�@IQ%��;>�U�I����7D*!�q�`�Q�5ݻ��s?(K��<j91������Jly�>d;�n2�˅��p.�5��|4u�1T�r���o�4�tK_�)G��Wc���*�bB�9�j�?~6߇�'�Q��~@x���hd'�kv��t�����-��ZZ�u"���D`&�q*:�i1T<��v����F�����@��u�U�:t�:���k�;��޽�V٥?���v��Ia�|w���$qg:���<���bn��<��}�<�)�Ȃ�/2@�1M1��)�I��y�b�PA�y�}*�U��c��/�z9�	�ea��g�P*�⅜Z�y�� ��$[yk�1:�>Z���T�S���4�캕!��DX����+R�J�I�-̒}"��5����S(�v�N���`I�����Esgo��+�נ;)%ه4��튦�:F�2��
} I	KͳՑ�|�X2��_���*ˈ./06��\����ʦM];�t�v�芳o�x�P��#g�{#�g��������7�3Xm)�,Ž��^Vݧ���z�_ȓ�ůqdi(�J��5\%/��X��r�֥����C
l��:vW���	v��0�/�Ƣc�4A�������|kD�߼��u>gP�����B�}R���l]�Z����`J�l(�Q���Uͱ���{9��$��n"RO�(��K�c��sg�r��xp/��7L!Tpr'-�?��0��X��8V�yJ�[�/����&�XR�=�%$*��/C�#8�B�.}D��:[�~}7tT���z�׈߿�Ũy����P}�< ��L�o>����!�5�{�� >�0~�	'I��I,��W���}�wCRs�ʬ�N�C��W�<�tU�$�;�|��2��}�y���D
�u0\#p��j�	�����w����@�Ȍ�����ҢD"�^^�T��LҤ��-i��P��n��1{���!��"P�$�]�̂L��x� (w�R���I~�`C J����G�_#i�K��S�[o�c��c�w%Jk�VL>�	W5o�:}��/�#Ǝ��M�n��yȔ�*�
ev�� V�w}��"�2��U"�N�7�~�f�/ڨ_��q��3R��GP�U"��o����!!��!��s��U��J�,�)f���%�ـ�tuǖ	���0<��HK�Iߓ�V�r1�T�+i�����u~�_��1y�v���V�>G�SF�GL8[۰�K�)��������S��T�F��F^E�+�q	��H�M��s�X�3�������I}�B�V����%�7�H��ݠ{�X�.:�'PuX dU���H�~�o�\�@M�֘BIvJ��ف��E��v.-���!hU�Yt�<�iF]o��NW�e������)��S���$m���mߩ�$U� [x�ᭃo��?S�A�jd1��݌;^���{[��_*�Hr��74��y���i���tt����R`h�i��*r�Vc�;Nq��i��A�'��`<g��n�v]��^������ἲ�A�B��?djNb���DZ:6Q��ƭ�7��
��zr}�tIl�m�s�>M�Z�%�����#V�x���x{{s�,L�`k9x��<�t�Kq4j��o�^�@}+�V��M:B����ġ�c����	�-��K3Qϭ�~��=�=�z��k��*�:��<�� |r_e���b�NO��|wAr�ЦE�|��4�8���>~���m~�'r��N��h��o���6���k��\�6�a���̂]ڠ�����b�3v�lE;&�u��n[e"�O��t��E�I^ oٹ��@��=o��B[�~��W�LF�R��a5!8)�������ι+�?�_��\�� B`�,Rrh��xŶ�����@�rn����;�����r�~��ֶ�� ��d��7�Vu��ךg�Wt��w�_����0\�Ḻr抆T�ͬ=H�q�F����@�[H�ۧ HF��pB��B1�P���G�PR0�>e�v��s��*���Y}Pp���&�'�R[�zS���B����A�v�*�����$�2F��*�v����e�ƒ޾`�#�T\Lѧ��Y8���Y����X���R�h��y/?ԑ�W�#@G���T������B��С�Ԅ�C�OM(���k�KCv�(41�0T��6K�a-�j�l4�M�75Z)y���)!Y���W	>�yX�N9i�����U��?��TK��"v<E��0��t%q�'ڭI��6��U6!||� �g~�I��S�ᳫ��]�_��oe���w?�;��z|�����Re�T��H�b�W4?�f�c����U��g��ΰ������q!s��cO����p�Ld'}�����'3��6(<�U��H�}�lU�v��fv������Mt#Dh�&U�hq����џ-,�on`�[:��G�J�1���-���8��!�m���%��ޙ��g��i��!�疊�Ue�V'}�S�/�pk^�}����[,��$�A���9���#<@�J��e4���m��� ��QÀ3PT�LȏG��ڕQ��ι���׬9�;S�3�l�T%��lc��<s��`�I�N�& %���h&�=tS������� k�H��cH�-V'KL��#�|��+w^צ(b��,��������$A�z��.�'`�ԝ�C)ߔl *a��_�ß5���k��� }�˦�
�k�ro�d�HՕZ�zG��%�e�6f�P>Rs��H�M���zs�m�u��u�W�n��@��6"�1��h�Oʭ��A�]T����A&�/�z����{�Qۊ�!F��"��d���+��B�H�霢Ud$��J��$�6�͂��U:��<63��ƝjU&�G�'�����o9��ۉ|���^���;�%�@�#�&B�dg��@*")M�j�E��'���̳GO�<@	�/�&A�)��ev����O��<0��#�.zm�Yzi|vq �'N��jPߝ�x&����J6��:���2N��뚞 e��Gr�Sp]�p�t�sK~�^�}q2�����x�x�6�U���T�Εsx��\���Δ�;#U�&=z_R���ӿoL^�'����\#�N5`���$�l�((s��.(	����!<������0V�>�X�[ueM�Ï� {�I�o��U0��Ӟ"5����9�($��,a�"��;ި���3G�� �`7��_-�
F�U#wg��zz�;������ �I��m���D-v76<�ߔ�������`���k��⏔����"E��b����<��˧����J�,ۜ�IO���Q�c+6E@k�R�qYB;wutR��T�� ߶��/���]g�H�����{,	4��m#����Q�4�7օ'U�C������0[��O����/��V�!s�jc��D��}���#�/��V�xr���dj��m��U��j �T�:t�@���h���UGj�S�
�oF6�=+@L���˄�I������A	^�k���j�[0ݶ�	9�*W��M��;"k����8��b~���^���ш_����TUj�ػ�0?�	���QA/�[W��J��{�Q;$�-0�;4��S���ƀz���zU�-ͥ��	��-E����U����(	�-�^�:�����v�eI9lҭ�o;�{���qְ�Dv 1�O@-��AA���\��B
s��#${�A���z��2s[`���Mg�L&��s/���B�F�wyC>8�?�Q^����hl�^ceB��B��v��+_`�G%��!��*"��9���8>�k������X����A~[.Xj�n_�V�ӈ��g�5�a�0'̠�$7��$�C��V[�%^.*�b@|��{��D�z���S1�w��I�<�<y��
���y���%B�6�6��-�)$��o��{�9�瓱�u�P� 2NᧄR�xe#1$��k�����b��� �th�G�Ow�4�ַ������p��s����IF���@~����L���.����!a�BL��)�!��V�D��1�M1�&{���D&)�O�p(	��E���0ZV�]��ErI�2���YM�K#x��2-fƀ���� p�����1
�?d��B�;>�O�1����h�W��o����)�.�k����Ng�eއ6{��W�_�v�0�鉱%�k������XϴMl��=W�H��R�)N���7w�ka2�eq��"��%	���t�jR���������h}0��nJ&3�	_�p�&�@�gG��1���j����=�p����g����g�\ʥ�S<7mq�lY{�O& ?�wzi�N�)ƙ���4"�;w:�t$�.7�Ap�F|�}��<-��Dn���j�oى�o	��-��������}{l���j*�6V��q�}PE�W�~��5�l>c�̶( j�d�Ԗ��l��gt��[��nԿݒ�����6��b9�:r������[���q��-!EV2sQ给�N.��?��Z���}�؋'�|F�R�6����j��MU�B���G:P�os����c���������	{��n����B�z���9�~^�l����z,��YeR����s�"wptKG��	�1dq�6�q�j�5��/�X���7���^ܤG�'�l����u����`5�wW[�9b�y�ᴬm�XW>�G�ڬ#�����e|�,���%�y>p�r��БggE��OoѮ���)6�Tv8x�Vw�n�xO/��/��K�{��cR�s��w�ß%|Q��{y��'u�����"��i�$|Y�ƪ���B�S�Ņ,�f��hoW�#�u��9� 8���|�V�G��D'g(��h��s�MԳղ-={s�ћ�A�C�^� ԧ7�y �[���־i�Iֹ5za`]-�.ʖ��[uݫ-�CE����נ�����P�H���Z""�V�4��
�����;�`�'Ik/����o��ij�neEӎ��������O�_�VRA����j���$�g�b;��Ɉ���xz�cCt.A�G�����/zp�3�m��a��ͭ#��o�'�z��������5���_��'�d�=,���k�����l�Ti�4�[��������Ճ�6 �y�k�Ed���b�P��w���;����L�ab���n���V�w��y�,[�A>��`;��n#m��E���GJ�S�A�[��j�lt����E��?�B��)�aۿ�R����߆ ,� >$��a3��8�+/��F���8�L,RT���^����*����p�����H�3���7�Gb%��n.�j���H�ebf�Y�CU�t�����T;#I"���2�������;�IT��9w�vf�w�H�rT�G�G�4����.7<F�e1H1D>�p�<p"����˟��&���ܸm�!�EZ��}�Ʈ�SЏ���DH�_�jY�=��^�%Wt�ةa���]R�t�Ts}>g�[�d9!EL �eV�$��~���K�o����+:o��e
��r�}ľ�7�lל�����zW���.������Ԕ� x�`@��WN-���/)�=�_�U%��'��x+�FWY�s0ö��������'M�PG�O5q�K4 �
X��c+v�i�*=�0ʹ� V��@��?��~�47�e�{|3�X��; NLِ��ۙ�LD'�31�e�0�;.JY�	�?���~& �W���������N��Xb�Bi���%o�ʨ ����������W�F#�����1�7~����s����qv��b�uG3oT�X�9�Z���N���>:��P;_)��*�W�y>.��#����_a>��.~8��9N�� ǔG���ꍏ|�-���4��Ae "�Q��\5P	����r'�NM"kU������ɇ���������Wq���ٚ��Ky%3�WQ8��Ua�CT9n��9[��JA�ChWS�tl�BG5����C_��]#��l��+��~�^�^	�JW�O�7��a��3-�X @�W\��NP�!"�İ�Ӿ(�����Qo�����el���6�Od��jA�2ƂM���L���_�L���6\ �Y�#`����9�Ǩ��*kn=Pɑ�:;�*��yJ�%0ծ'c�a�,Ģ��\d�e�Z��p]�����;�c��Ԁ/��D0�}�>�%x���A���R���%������{��#�P�Vh�+�<|˨+�t-ªmD�X#�X�Y8pրT�3�`�uy���{8C�X\�["%]��*��B�D��Z����I�J'���8�'0%��H]4�Ġ/��P%$�WnI�B��JSGi��*v�� ���:n�C���qH�^����P��FYa��	,���x,�����z�S��P-��OH���QG�m��5���`�� ����Z~Rx��2^�p�6X��6����gX�D���X�+�0�:H������T؈u����{	@{4�ўCy	�X���v��,�)Ck8�M��/L)`@�d�C��ѱ�Q1Ҿ�LǿC�,���gQ��K�>�|���l��y;n��[ �A�%�����A'_,h���sC,���&������]a{u�8�ӊ!HB�Va���C�1�$s��y۠�2�/��5��YM]1'�r� vu�Y�<g{��Q���61�87ߌHYۺ�8sv;Uk���7�~���zX咃�\C��m��ɐ&
,,0�"�z��|P��F���G��Ҫ�q��c�G���N�~���]/���p��ۉ���5��p<^��1@�(�m�r�rl�#\jW�G�1N:\���^@���-���P�A��8^S��/w��M4�z�12��q@��}r��*u�Z�P�C"��{&̱�ǳ&�:S-�"V����#p�\����0��=78���������B�o$�%��
���;�})rA�x�:�����G��X��I�+��?��|XX�_�X?ֆ�Vd��Ao��4`����E�G�7U��٪���6�窯��28 �W#�tU���Z�Y�;=PEy��2�y�� ����Z�:��t�9��>~� � r��� �|�H-MC��u���|�OH�G�}�TD.��@���B��w�*�-�zl�SyJ����KA�G�����R8�4���H�[�KjQ0[#��SG��S��p�\�A\�֡ѩ_�����m ��W��x��<)��+�k#6;�����(�V��t�(��}?�S\��!PNNo�xd��}��>fG���fJ7��b}s�xu�;��z\��M�=��J%[�<Y"�ޑ�b�6F�N��qS[*J�a�A�A��Ni������}}0	 4:�Rv���G� �R�z�y0W�3�C#w��FmN��]P��r�)k!*�\�r�MYa��Nw0��n���x��8�ǨT��M`(�F�c�\WE��Z�-�o�}�`4!9����I��3� �p;}I3�+�6=%J��3�e�IF��d7�Lr̟$
	��I:����
�@؇<K�'�{�;t5�
�4�*�d����-'Os������g��=��$�����5����n�i��s�Fo᫺k�ɸ���wD9Wڐ*⹥Y�T
w� ��d�-��\�"�����O!H੅ܟ>�BV������.����r��R[:��~��S��a�l2>3��x�F�O]���%���l���?���^A%M�A��Rx����c�y��P�;�G�N�XY�D�q�@�f�"^�[�ۭ�Ѩ4�L�w� �����!��ͭ!	�2�3�1�n+��L����oh�3�)�*E ��\�aܬ�f8w��RT�4��͕�R]8z5�V̽��5�!��:��F��g�СQ�kH%����jp�\�w�8�"W|ք�MX�{��3��Ё(*ߙDC�i*��!�}�S��A�_�g�^�J�?z�eSP��/]X�>����b��aF&�Z�2Y���6��d��e��f7%�_�ܒ3�����,��&�ö$X��7)��������Eߘ
U83q�^&Ğ��b��
k��̚���4��X�{Ap�������T����d��̼�%<J�Y�e�0,���] HM3��~�KFh�>���,@�\����5�RH
L��V,����.W����� ���)�R �/�0�,z�%��ِc�wo�*K�簦N�����i��`�]�>h^^'3+�I��U��u����Lr��~%�������f�Kk�LD�SPR^�k�'�W��-Q�IxjM#5��A�i*Sx<e���[ȟ��Ί=T�,�1߈jd�Q~��;#�ړ��.zGd�_��ڐ&�0���O�q��П�޶��W�o�zf�f�}Y�OI�]�7�@��r��$P��]���6�K� 0 �:���� c�,d�����t��#�9�� n=���kk����]O0�d�-Rփo�U���-Ȩ��-^A���m/}:�=��>s��_�t�JH߈���e'��J�g(Ԛ����FNؖ�Z��q�����Lw������