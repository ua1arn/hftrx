��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p���d�������C�zT]�iK��
�@<�ю������|�U�o�1�;R����I����BSO�|�f���;�oά5x�,��Rіu<����b���I\���(rRׅ�O*�S���߯�����!����v��~f�s\���2~�ԾY+}?Q�B�9�68���Z���{u� �&��X��e���P�����n�
��s�xYZ��GX�GTaj���s-��+)_��6g�ڕC�������Q�~&燂����j�+F�B�A�O3ϣ�Z������[�Y������V;�����������$��0�?
�!]#�︟u��D.#Fm��y��ę���G���"ը?-qD��d���h���ُr}���||���
\�Q 2M}�H�)+9oMփ�{p�V�
�҄�Vm '$�_���@�Q�E��p���Z�W@��V���}Ke�� ��g��~/�����Q+�MI~�����.�!�OעKK���NM��fv����S��A�'�g��x٤�d�Iͥ,o�n���Eک04Ք{��.![�MA�e��
���^i�- ��z�����E8͆!��z�*Wٍn֠?�cƗ���NR��>�)�u�̽T/�-�5Ԓ^�3oh\-�7��< ��?���t�mf:E[�U��}��"C��,8�W��3�cg���|&�6�����}�]��i5�C�#�zR�<Z� �adˮE"��M	y����#�d�y{�<�-�����ouR��^4ӽ���\��=����aK���ߛ>�����vaX�����$rSB�[��+��N���.����(��?�]����oԑ���P�Z�5Uzia7{$��˃�rX�3��B�2�)�RΎX�ʀrO'��H�z M�	�G�>㪂��d2Q&�V�rM��*t�n���D�����FAz�'�'i������}g��PP�|�.CW	�Oi��?3�o�����b=#�-�P�H7se���Q�: K>Sg�nX��3H ��].]��#վ9�F���7��g�c���I�ҫ�B�����!<���Q|Ȩ�ͺ{�!B��E�����w���y��AA�"�5;�HI�o����Z��Y�B<���{�-_���rVG��qc�%l���Y��"��%.ߤ��M|��t��ɾ�^���y �C7�5�M�_R��B,�@�������N~i��x"���B�O6���������Ա� �@?@��kk���8jn��f.4��2�XR�n1��^FVA2��Jٿ����e���'�)S�mhCd@��ށ(�����.h�������������!����q�xX�+]v�5���䛛�1Qm@��	��o��[���\�-A�'+v3�y��n���6��&�M�[�"��h?H�H���N��z�Vyl�&w���LPXA7t�[����o���ʆ�N�Y�b	wɖ���"�}
3;��7d��mR=����0�r~ģ[%l�~�Z�1#tl����?q�&�͠�)w�6