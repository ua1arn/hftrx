��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K���e���c5�B�s3!S��s\:=][�*��7���ƃ!K�Q���ݠ��۲}ͩ�<�>��>+�J��ph�m@ҧC���9*/�5���2]R��L3�(��}����0�$��O�-���"8E����c;!L��x���|G�F-�3k��C�����#WAe5]o�]>�G	���"��&3�*�l0X�<t&��;�G@R�AB�3�����[3�8?6�SKm�,�b������m����?u�����Y�����ppf;Pb@��w7�%O�"��.��$J'��2D��ּ[�Z�v~ЂL��[��sx^����a�Y�T�5��d	�|(�=춒šH#�)X�6;^�7�����"�V�c?��rc��!�����p�8p��5P�&ᵤ�Z���l�z6_��[0�1���}i�L�	�d��F[��W��c3�P�N�r��R�~��E�w|�J��p$����o���?��oDf�õ�X��<r�3��2�T܄�[�6���̽�U���f��w�3h"�������`(P��ݐ���@6ad:��*��g~T��R���"LFA���t�ě}P▍�l�S��� (�y�UHP���V�Xٜ�̈`o�=[�W�%���q�H��� *w������r4����y�S0�mQfAb�2�:
 iT̶=Մ�uP,�ʙ��u~hp�0�Sxo�OX�^X���d燢�5���X�H��2sa5ԂI;2��r�7�5Β�wg��j�&IW��� ��d�({gZo���d�tUJ-os�W�|n���1��G2�7:*2Ē��Xf��ءע{)�
��ZXa���X\d�_.�]� I�{]�����!s���mw��b�n.V����F���ĆL+�AG�kCQ�<��Uh����ab���ȵ�`LE��*�����q�FR������[f�uOY�6� �)f�D}h�Sg�a�M���7�q�	w�w��}������:>�!��M$K�h�L�o��U�;���̬�&}�)�ݼӊ���{p\�����m�\{0� m*�3rQ�%�5o��:��r$�ls��Bsd$3���:��c�X��m|�eM=\�j)kL���!,�N����t����z[/���a
D�u'����A.?��lNR�&9
4Ұ�NEY�.E'��k��<����6�G�y��=�}[::ՙ��uq5<d���{���n���
���=P)��ys*L�ċ�A���d0�(����k���_i�Xo�R�oY��U� A����>#v%�3��� s�
�r	ta���܀���R.|��w;{��ۑ����T���h/i�Işoe��7B4��p���?h�������������,�4���;�{Qh���+ܝ_i|j�/ ��]6U�+-a��l��V�f\�kz�1��y@MN�:r��,y iÔ��$��)�}_ZZ8���ם��=����n�P�j����l����Zd��l�����l��T/f�(����xDg���/��廨�ѓ���Ih<��9D��}GМ�N�Gxu߆�qU�NZ��(��As���6�2�
l�b<�n��!�CR��'t^�i1!��5�̵Gt؆��S���-`ʋ&S5mIT9$�a~�-;$.����i�"Ta�����tV'���X>?�����{_����vy�/ c1�K�C����Jz>w��)�<DQ}@���D�-_&ލ�`�\����������]�M2T��oq=�[�p7��	�7C��)R� 	n~-f��@3�t�P;R>	"���Z�0�N�_0����n�r�O%'�0�>g]�!��l��D8�;�R4��*�	awUx�%T�3*s�q9 >����!r�G���/��s��BžG���P쓭G�dN�C50��N��{P��b)��C�q����75 ψaU<�q�䴻1�v<.#��>��:�NBbkV��c@/�N�����=��],���Dm�Q��׋)�6�g�r/a����a��d�v���JT9C%	����A��h�X��d�I�j] ��u�rd����������1w�(�rd�j���kM��1�������.��1d_�Kl�1W���8g벟�S������#��G�����Ep>��9D_$�1i���y�Y��.���Y�ؙ��&���	e@�KU5N�7s��J��fJ#����� E"x �Y{ad��Y���f�~ft�1No?����P��(m��� ��`况"��@��E<d����~	��i�Eu�O��Q #E���è��θ{�=�=[���aU	��+�@J�q�=��`9rq��k�&لu��6�0�]��/!�bo�Tɪ����d���=�k����mp�2嚑n������{_f�3�j��r�N4�|�iX���F&i��J�^�{ŗ��Qk��5�.��ꇹe�<\����<J٨x7�2{݄��)����̛bN���"�^� &v�m�L��\ϲ���~"��A�H|L@�ѓ����������t��w!}�N�b>8�e����#���Ҁh�	��g<�5��P��ۗ��5�Od_��{!R.i�W��h����h;.�"\��ėI������cҪ�� ���2�R�x�K�$�)���}rd����L���)��G׵�QK̀�gv�c��(
<�"��Y@�;+>�4|�
���
s����۔��F�X��	�hve���Ȃ鵵t��@m����*㉼�������x,�|��Z�u���v���Z>�'�2P�@���wZ��bYFZ$�����<���Oj���p�Z��E��+gle���T���p��W����T��j�BdPDI�%�Ҷ�Lu
�2n{�""_�(�6.V���L��8�k�������4��jD냌����`A�uJ�eI��H3���y8h�$5u�>�jq(Rd��{�(_��Z��2��K�%Žop��I7�����a�#<���� ����Ǖ���K?SѡR~l�?H�CaEJ֔0Ŋ��e����&ll����.�wE�~�Cd0<�~���N�i,&�a�6�����,<A��,/���O;��� �5�+�V�
+w۟����^W�2.��s~y8$���_O"5��/��R(ru�#����4�E���?�~�BC]�I3\h���\�O�DBȐ��ILӊ��)%�ܵMLػ'H��|K8���$U���a�7)J �W�/o�������K�����7_�? {jM���?�]D-l�� i���A_�8�Ez�`(fP����!ʑ9L���� �ُ-�)���3oG�������&��Vy��m_W�ο�����Z�� .h|�rj����P��Tq��p�����ά�<����_Ճ��.8K�
������0��%Y�����Zw�7~�v�K+�Mj/}��?F�e��O�!,VƼ�@��@�`&�{j������B&#w����x��n�ጆ�5��B����Zf�G�=ӟ�p�_$�>�{�Me�%�w�>Y'KK��S-YZ��r�>��K�jq�g�N�ɖ��P{�,�ʹ��憃���xd����<Im�^c���EEOU�9=��a%�5�AA�n�W2M�{��-�dB-1?�RkZF&�ǤA�C����AF� �O�y��.�|r\�E�c���]X�m�0Q>e����*b̈́�>�e������ D��������m6?bɝf�WT��0.�o����?_	`?]�j�?Y�Q�-�9���_���� ��
@%�g-�����G6��Ӗ4Y�H�4�<B_m�崲�e���I��n;B���(���UVh�F)�v����W�8���>��O%�hێ�U���$ݶ�؝�Ъ�|F�� 4б�9߇��Xݮ�v-��u�c؝��k^�.{6*1:\s�^�  F���_<�\m�S�/��͡�t7W�-+q�>-��Z҇����x�Q膼B�kǰn|E�0a��"F��=��<l��^�*��|C�A�3u���'�_��Q��������hutN�ݐ̵���Nb�B�1,q�<���������`�܈���J�W�C�	�n���e��x�Q?F�i�P��[O�xh߅pA;��͓D�7��@�a�QX�L�f�TX<Є�k`��ط��!^c�#`|��ܨKҋƹ��>Ft�� e�N��j}ԕ�&�#� ���}.����Ɏ�m�hB1&�X���rd�@+X�_D���;���;�<I��mmi?��nwհ��Gч�P�8~��{�.��j�Qv��"�_qh�kȾ��`N	)���qr��tX���ϝ�!�*�N(�7�x�5=��e�Ƞ�fڗ����7&D�w-�)[L�m=�r:r�w�.�H�q�"��y�l�� �c��x���0��J���6�$���Y���2c���aA}8��V(�c���h
pW��|.(O���J�iǴA�*9��9�X�W�~X3��'��%��Ы��~�5R�y��!���L�����z�����Rk�T�v&�oMYĲȭU�xX#�]"� }��a2�l���'���L>�<��I��`y.f�*1<��Ԉ� �^3n��t��]��T�6V+!����]e�E��m��9i�c��:�4�R��J��"�����M�#�K^�l�`���54LBX�����j���z�9�nb��T�a�W�L�~��A�g<瀸�4��I���l��1�WFg�/�G�'7S�� 0rpK��`�4�u�P}��i���ܤT��t�����/�!���OH_�VB\I�����T"�fѡB�'ܩpr�O�݀lw���@>p~~�E�i1*���
���v�1����21����to�E����n1q�?��\�����WQ�N�b�ߟ� ;�u�w���l:f�Ҍ]{��|�uA�Ecڲ}*���vL	^ZUX���\�&��C[�Rm?0ܴ��޽�����o�t�gZ�8�6�%}L}8TX��p��Ͱ�":��s��t3w =G�G����>���m�J�c��n�	�[j���հ>���d�H���"5��䊨T���v	�.)�m��}gY}ө��)px��at�#�X#�\aB(�b	ֈ�5����ٮ��mg�S�IE�b� �޷����O������_��;h9����
.�����pANk����l�pLXI���MD��ئ���jm��w2��L9pi��A-�)��t�Z�����
� G�xWV�[�Kj�SnA�;E��uFR}3�1evԘ'���f���:E/�;�|{99����=+�5R�-Psw��@��1���t;�q<.��%�i9�����m�=>�V�,��W���Dd�ž-��y�Ӝ�+��飩L
�V�%�aH �ԋ���t2@("хFs��4R�O��t�HӘ���y��:�Z������O�d֟R�/����l	Ac��ڤ�bY�n��; g3;x�'˴��w�҇�!�X����gl��#��+��*�?M^�M�c�xc�C~@��e��v�E�M<x�&@��C24�8��TԾ�7{~}e�R3K��Ӧ��uj��
��c\�B��?���=y\����6Q�C_oJPb�	��a.N�g��/�`2�MI���`�@3j��2{��]t'a�N��]-kϹ�u��e���;�����z�)�Zi��fk:���A����`�iV�7*~���x��9�A����'s�
)"<P�6�E���jcL)�tuo h۪��d-4�8|\�Tnq����7��ڠ���k��_f����(1c6C�d�V�̘1�ikێ���3����{4����rK�n����{����C�KD��[i����31��m���}�>��� �S�� �^ُ[�9��@3i�1��<��^Zy�UX��%��v[ۧ��Af�pK�ʟ(͹
;��0��&�At��l�	^��冗�B0w�k"�|hx�ĮJ�J�w��\K�P^Ĺ%�L�z`�L˦^cz�����ih�����֕}vVs|R�`ag���F�k<�;��C�vb�
�$
����Y�������r��Ҏmv�	`8�p�M}�3O{��	�V�
S�
�V@�n�g�w�$VD�?�M`v��*�� ���2�=�,mt�1��a0�hM�4��]G_I3����}RmB�[Ţ�3����$/��J`�~k\�ĉm@ �`P��tg������>"��}5`;,��5�IV���j �&˫�o퍁���A��M�˯۪o�O�8D���`�Hi���2q�����& ��պz����࿎,~�!n`�{yF7���$@�1��O�`���Pt��Հ<6~��Y�ڎl��������T}���u���G�'A�N�	Ϸj#�#���K�B, ͷ_ԋ>#V����h�a )���N9ZGY�w��3/�Ɣ��:6�K6%�/�m�`�#��������O��a�l.�Q9�Ù��e�r�q�f�ځ֠h�"���"��'�z�j�g�)�&\:��*V��(�f:�ard��5M�T����cXY./č�֥5�?N���=���Gi����'�JnI�B��X^�=���s�J�ijq��Z}�B]����ԭ���].\V������!��+�ĳ�"YH�P=�>O�窩�NWH��n6���[%5��(������u��bl>m|N,�VR���2���M�����xʈ�: ��M��zD}��Z4�\��%�4�-�ٳZ���^K�y~��>ʛ��yݬ��]u܍ԭ�����5BDZ��o�P����D�qAV}2D���/|�M��,ގ�Ջ�3���Am>��zV8&�i�Fk��|gY��IQ��$t�R��so�^��S��;�"F�9Q5��"a^���-�G�u��H�v��� �pT�]������K��g�r^A6�9�j,WDǦ��jV���>�q�ꌾͶuStX5tZ�l���df�0s���k��Mø��g%_e�hH3PYD��6$�P{ x��6�-�wYS�n�J�CN�]�b�)c'"'�!o;��LV�1-VDr��CJ���I�K�7�l#�sv�%l�|��s8�0"!d���i��#�#~@ůt�i� ��j�Y�K��+2�6ĩ�}�	q�Db����>�KZ�P�BLngsf�^��E�Boн�����e P��������p�.���9:�� O��Ȃ+��F,�\��ѦZݮ<bN�����[�ơ�X��n��	W=�0�:����Ro��K����}h����X�y�t�GZ'��l�5n�ԣ�:fxd��h�I�ݗb~7ύ�1g�;���J�K�2c�\(G���������o��#GX\�,pPI��Ė�D-�T�е�Qחr�SuA���*�%�aBN5U��2�|����Ͽd����_jV���p��;����1�V��r`�SzR����i�2��nA�X=%�2�'Gռr��7�E�%���ŏ�!��U+�!��oo��V�ݘՁ$%6^�Gz9o�[.B��"xV�~� tc���9��QS}y����j�ya�LP�R����Ldd1�3���T�����$voo�E���^������9օ�S:��>3-�w9�$�+-n$q\�3�Ӌ2�I�RPYPQe԰�Q������|��'�Y��[yn�E�]q��w2��αp�'�������$��"�C��k=��r��;�|��_�!#��-x��g�ܬ�P5� ұR�K����v��-�#y��%ί��"��jF)�7�9V/�8�7v5����7��n_�1,��&�i��n-�'�gy���/�� -Ԃ��l����s42M%V�ŝ�@�I5x"s�����6G���~�4���N�9Y��<	����_�#Q��q�!���u����;A�'� imFne]�!���1v ډ����䮎ٻN)�Ni�*zkuS����(�(i
�*%�EFvC��'��+��jV���o���쮐˔f3!��tG�����x��XE�z69l˜�y�>�#�
��#�]�{Q{E�����ͩ�Wמ��/�nP���[�NFd�f.=i��p�}�eEF��n����r��N~�~o: >d��I���h�s�䰺��L�
�����n2�߳�/�0ן���~�X�\�[�ZL_i���׫q��j�^<����|���"�ϸ�:��F���l,R�uh�{Gn�]��p4��ɜ���,z�W%�����ہ DS#	�7��C�MC��C�OQI��C��(�����R� ���t�oƅoT0�����\���������Ί� f�P𢡊����>�Vp@^b]8F����[K3uTf�ggO��${H��;�m��p�<b���{������섣[ȿ50ۋ)0M���g�U�h: �@�.�V^AT�+�栭�=1�K��;.e9�|�^Zk�?ggTB�Ă����"�HM�xbP��`<��;3>;T�9n>8��s�SXύ�}ϟji2���R%jHCm�o{	�]��K�}-�Z�Pq��2Kg��U m�4 ی�`%+���p�����j��r�+�tD�[{���[$���03��pǍ�z��
��fh*��/��Ia�J��\�u@�S�؟?��xI p�O�.�҆5��
H�,�����h����3��W�;?�xQ�0a?̓����/�Mp�� )�M���>�@A����g���=����>�6�E������g�1�t��
��.� � �&�?�j`H5�.T8�+e�J�|+w4�UK곩w��U#M�{��9�[f@��2<���udI��u�w�;�C㏺����[���$kKw��x��C�:g�4<� �9~���k�S�������.���8NMMh`�0����*z2?}�6X�J!@�~�]���c(���F���@�ݗ;��4l��咠��#V�XvV\K~?]n^�%5�W�OË��~�N7͈�Y��SO�%q+�ڎ�ɛem���(���&��XK%I��5 ��&r���OG���%&�6�<=C��Ѳ����򛳵�Iq�L��iq����E���5���?F��rB�B&��g扷����V�Ӱ%x�Y���**T�A���r0�G���'o�W(xȮp�T�)���F�_��]8Ɋ�~��Bl�4��i%��4]6o�"/��6�߲�?5�I�cۄ�Rl\����3}�9h9��N1~z����pG=����-�����L(���>�c��i}]$�S���	��6'��,��^0��`LwX�B�T+f%CESp�0�*,�bsʎ¸9���Md`R���&mF�y�gL ��ò�0�����˘��M,¾b+~�82��O��e+?�Ezs���F5�	��g��]�� ��z��󪎒K����-�\Y��b~Nf�tRcKlJȠn5%�%�1�$�9���ʰ�
��e,K֖�,��T��n��%�G��	��|N�1_|�Wc������ĝ����!�`��N��3�>��VQ�s����L�60ŁR��aK�>�H2���>Cmq��!2�q��>�>�R��F�8A����K?g�{�����I#+�Τ&��k'2%�W�<�������PA2�e��Gs/		�9m�j/�zq�`�X������ �������d��E��3<������r�6T"����S%F�u�}3��O��5X�!�
蘢�x��<\�S_f�������I���ȟ=��~�/�X�'E�f�t�Ex/pV�J3���;o e��?�F6�����������x�S����eV]��M��z�k�[�Ӈ���6gO�l�
�UR�k	�`��]�R�Cc���+��J�0��}o_kwܜ}��(*��t��$m3$��Y�Ε�6@ھ0�����i�d���]�(B�m���@a��hB�X2��x=Y?�h���=k�����ӿ����(R�֨W�$�9D���,�9��Jx٤;�,�"�&8����l�7q6����P���_��T�����K���:=&'�ԻC���Kml5���~��2��� 3�I�jm�%��K-�O�o>w}�,&M��E�Q!�7�1���T�8�����N����P������������h�(�۴=��Ϸ@'b첞���^"��|X����tN\vs���B�
�g� �F	f���?~��=�j���"��b�LO�ΐ���YM�����R"S?�'��1Ά�p��T�W����F6�m���U�9�������^�������� F`�B�7�%�M^SUC��e����K��c��c�J v���r��[�j�(  ��
���ؿkȠD�+q�}���I��a��䪥�f�M�EoJ�P�c��o���ݏ;����\H�n�a�x�&�g��O��e���рN'��R��3���V�"�3/H1�1z��`�ld_5W��SsUnb��C}���=H�i��nm��m��$���=D�E����7ܿ6��j�U��WA�풨�.�d�Hrv�7�~D]϶Y���9e���_u�Gi���?�<�:�����-ٖ�\f���AciO��x�G��f�L�M�m��?��,Gv{,^E_����9"��sR����5�ٱ�L�_z�֑�y��k�a����6S��}to��d�L�t�t�J4����~s�٪2\a�_�eX��F��m,p��C�)��z%6�G�F3#�C��Z/��0�� ʅ���6�C�F{xn����t��c��GT��A(���^ך'#M@�� "ꭊZO�I9p*�nn�2�JL�䤆?���\*��6�T=��]՛�9�o�%^�����5~F$ߚ����\e��<��)�=k�Ё��GX(�^��x��i�X�R��r7�u�<���(~�y�+�@g�ޘػ3J�6W.��1
%�P���I�4:ɿ.�Zg�����>|��~E��:�J�E1�����<��SB1@�Gs�}� \D�"����b�ma�\�=%,{2I6��h:�����,�uLl���Qq^�7�
��؏�����N�0c����v�d%O��k=��.Mt��;]߶��/v�$L��?7�,�J�����HT"C�:���Ve�.fkr^��,�ە�+��IF��ֶH�c^�T��^�� ��H�����X���"�	R�t���ңS/�5�J�)Ы$9��ִ�5�c���އE��~�%��YR�DQi�+����Ĩ���A��Y,�=��>Z>����u�A��	K�4���I6t*5i�U>�q���l�v��τm�&�Lܛጡ����a��