��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b��%[��$~�LK�x�c]'�Cj�i�7����$#��n�#�@�)(>C�)ͱkႢ�HE�U?�/v�j��[�$��?�㠇˟EjC����>��]/E�;�e>���s(�S;���)՚�o�D�<�F�_`Sq?�`i�AhKO��#��_.���zyl���v�dl�K��}���Q�ao� �2�О����þ���?=g|�E���ʓgϨ��9A�<6�l�l�x��X�_pY�+�]����{��]"����ik?��i‴�	�{��aa�^
*I��Î)�3��JF����U�<$�G��dk��	����Ǚ�����<�҃���x3!ϙo�q���}\�&j#����l�E%�Ԅ0��}����B=�;an�Q�@BO��~�b�]uÿݝ���|�jw�.2��G�aˁ:Y.j��1e���	�������;�@����\x��V5�aE���_#8���-�#dv�6k,q��"�!�;l��@z�E����A�!%ӽ��:�<:�,xC�)q��&q���f�Z����?��W�."�+�}����΋%Ё�Xd�6�u����@+���H�\U��!o%R?�kwTm6u\v�/��D����z���u�"�3����U����Z-��%�Z>�N)��Q�K,ќ�\�I�ݹ��S¯�ؓ}� ���n�Y��tjI��3yHZ1\Jr,rf(�W�.��٨I_Q�"l�r���
�2�?���"�h�]�Ą*��Ȍ	;�Fz���ni�Pdd�c��I[2~c��F$u�������m����]��r!w��WcI�N#f m��B�#[}����Ub��h9v���	�� Ň��2���q}�*u~���Gɧ5���'�
FgoX�82�k�]�"~��)xl��A�8�/RPa����*��C��?T�`>�S>���6�IֺS`4k�F�I���#iE�]K��<�`��b÷Ϳ�A�6�6:c��x�ϦgkF7l]��ĉC�r�����{*����?Y:T4��d����A;u��ָ��f��1��<K~�9|���,$}�3��y�CF^7�S�a��J�d�[-��;[�6�tϾ�=�/�"�,Pf
����������
���@c��7���y�n�\2��f5�-xG�,�0�jr���8;f�)�
<CV�3����E��6��MQ�&�ۀIp�[�����3D��mYV��U<\�掺\	dV��ٔ��ؽ�R��F�me�&�Ǫ�/gLuǃ��J�v
��t
m��F�����`�������-8F�M,.�#�E�m���M�֧���
n�;meu���F,]��Yʠ<�}'/�/���Kg�������RA�W:5'FO�U�.MYVgL�<�ݙ���>%��Ȩt�N��=o�)���**^�F�1�G�����W�UՑ}'Iy.�̙ڏ��1�g�����J�~sP�4�º�R�*?!';;ߤ�{��8PȦ��t=$}�����'����p����MՒ���0j�ά�/��ږa6����LaJ�q���Ë�3���xġ��7��/�{L�ȕ�`�G��s���\��=�	����K�V%R��{t :C�a�h�!�N������TRC��1AT$L���!�:m̫3�|�;�y�O#f��h7L͸5.��f��T�W�k������Āк�O�
W�UM8�JՌ?*���`|��� B�������8��� 0�.:ԕ��1��3����=�.쇕��.���V4p�Ϊ+�
C����<>}&
�9.��<��/_�����k�0a9r`%�H�"���pAq��y���?Ȭ��욫ٞ+�AHћT��P��Ӂ�6�<o X��2��Ct�9La1����A|j����9�u����y癢Z�%�7ACE	i�\�n�s~��y��n>Z�� ��,�(�3��>���q<v���19&�]~K��k��F�S���RK( 6 *��s�;DJp��nDh�hpp9�]��H�C��w�<n�	D�i�MQ��FDI#[�U�ڠ-�����5�b�`.�Kg1L�0PT�~GvUk�����ް���mI
RtTYX���j�)�4y�����G �`'�@��������tJ![�
k�;��K���)d��9��$���}�����lUS>��[���n��r���+�m��PBO}�E�%��tm�Y�᧤>g���=�y-��S0���5�n�ҩ�������p�>p+88�{��|P�Q�S�%�IO�x��8���:�����1J�j�&K��I���F�\�ܓ�jf�<M�5:!�pU��T�q�w�u��bc��F����{�H�5�f���#~���O$�������^�tk@fk�az=�݌���"��+�TD�
�&��P
@Ǿ23ڎ��E��9'���3[���8�wfT1�|MG�V�ښE�X-�$�s�� �H����o���]���:6�&�	��m٣ZX���
N�c�f���N��s����.ۉ�,��?S�w�j�'�8���Dn�&(};��\�	�C<�7���E�o���?y}%����{�
 �Im�4I;�/L��L]n�~O>�|�&�+�%P9�G=�իTM����C�=���L��_�-9��#_����9 � (��)�Ӥ�Q#�驓���O�[J Y��À������ĺQ�4�S��t���p�0�����q8�p͎͂{Ӗ���c�����4h�N߁%����炇��k4��$"��q-��8h�E�����/��U���~�=A!_�DeՎYڙ����5���:9������g�{[r B�1��b��?���}6����$�1%�X��Q���,w/��K�XF��'�
�νW��c�tc!�� V���I_LBDD�qq����_��DN�&������ �}�dOK,�����$rJț��J7�m��7�G�F��~p3��x��<�1g�/"�c��VJ<٠b��܇o=$��N�c��]s�d�;��Nᣣ}��jwO˳�T0��"/<u@�Zhi͸�vO�f	�����|̌�a7��@��_Qˌ}lQ ��lhK��L_�lT0�j�=3�kU�7:�uAL@��Q"�K�d��lQ���Y��m���iaU��w����O�;;�.��r�l�d_fh��q�ȼ��g�V��j+O'��9hSj��g�/%����!Э0E"j�����mU����edX�_���ye�/�%�	ic}�[��d[���=������u��OD�]	U����vAO�"XT�1`����g1�GXj�J]��B`�"�)5�f������c����\���Ձ�6��̼���MI��|tQ��^��.�@�S7zsTg"|�OiBv?��2:�p��p�E�O�׺s�� ,�1xs�8������Wm)�C��}0޸wF���Ǟ�E�:��v�,�7�%�=1j�*��Yb�oU�)-Q�5�Z���[�u�&��H8�Ai�4	L��$U�-P�׳�߬G��[u�%��r�0�'����h¤R_n�iK��7T�KH�Dm��oI^��	��L���_'��paL��Iu�2�^���#G���3�7�Pj�и�O*�|)[����7)tK��2��aV�@�ŮE/��+�O�JW��	�+u>�ʻ�5�2}��>�����ଈ��Q��,/�2�Y^����)>�<��KX�c'��m����ى1�*+�4�� �:��20j2�������:�y1�zB�;�E���8���^��~��!���P��֓Np_@z�ڋ�l/C��/�Z��jB_��,DHi/�k���"�� ]�Q�ڲk�_��$ו7n4�CXL)�΋)�}���A�.<���هx��&��_�j�"��)Zͽ)P9��$/b�(@��K�/�(bW[��~BZ����&{�x���珠��@��DU�f���-*�������`��_U�4�1&7ӊ�ݳeJ�z<Pnw���@)� )��[;���xg���*+eO��7��x4,�u&X|�#}��`Ym�=�|$v�Ѣ
���B�<_k��������� 9(FS���L���Z5��x����ޣ[�]!�:�>��Rn�"�_���X��riz��:�Ɛ}Z�_����ʽ��61@ۿ��,��NT�2�I��'H�����5�ؿ���!W�3�fAj0i�k94~�^��.���s�O8מu1>�k�O���dVs/"��=��&��ty{�\Κ���"jmq�F�k6t[QDokVD# <+L*'h4кW%h�L8b�R.�[�l����Mu� �D�i��1FGwse$P~b�8Z��n��D`p&��k��������$���[�O���q�ӓ	G�Y�	�ܱ��8��Hp<f=d2���$�}ʗpP��:�%���ҕ�̿��X�8�ҳ.xn��\��ܬ��5'&BZ�+sOM��#Ѻ[pR�JF�EAx�	��=�����P� �aQY�d!B1��r4�E!^q=+93�_8S���-1H#eG��3�!��Нi��Peղ`���XN���>��0��1����+��y)���^�q���7iP����`t=��� s���Q\|�EZ��� ���<��daq�^�mxQ^�/�h��]��`<���Ӫ3��6����y^ M�l�>N�\ ��@}[n!�|e����Gn�Oȵ��w�Q�'�cVx�y"JD�iME�ײַ�|�U�K聓5Rϐ�YB41��Tct0������h����[{��U9.M�V�������Y���_h6(�-p�~�Q��U�P�=�����Zc�	�g�̚�k/��Hz�����E�G,(\q�=1\�pgݪmB�e�soں� ��G���"f�s�Wv9j�6�q?������^?�.���A�Z��.@�$�'�ƒ�T:�ȧ���x�Z������ປ>�q8ӻP��������v��S�2S�&����z��t��#��n�)�ޑ5#��zW[� Z�%���xeR<�͜H�A�*)�a��B:��v[-�_�"��iNC�"|�zQ�ۅ�u_\�����s\��^P���>u�uk�Q�-XI��y&����أ�|�d��kJ�7��=�8{㻬:���D���lPP�A���~��1�
R!a8�8�1�f�
�')��𾧅�a��n0V�- ��X�Ƽ��x����0��!��%�#�r�д+�@Nw"��K�ު��%�'sӺ��KQVdN�Ȏ�mo��3'S!��p�i�B���2.4\�
���[eɋ<R�}��*Ϝ�6�Ӈ���I�]�+.��l�djHm��8���+�O����*)��9&v��S��h�c��q����)]dKnE�Ձ�櫾uU�9ܔ�̧#���P���&��ˑ��a�`�|*����>�Uӄ=c�7ֽ���n�<n���g��3�L㡐���}���u9;B�+l��¬wKG�}�_����W�	`=���?��o�QVl8�6X����-�+��� ���K����It5m7P����yYpGm����_]�AT�sޗ�7;�FX���K��IC���y5����U@�9�!e]�q&���Y�8�}�{2D���1W����h������,&z�/�m#~g��b��H�&�z��fכ��LZ=N\/A�r�"���������A����(��%6�vL�T��Rd�-�ѿgQh�����/]a����v(w���l8L������}(毴�f�G^�f�A�d)H3���T'��P��p�K�֕w��_���ءj1N.��g#��"����y�\����?�}{iT1
Z�g�J��64��fB����������*���鱜k�=
�p�����/"B��]RB�n���7�|��i�_[2R��uNwg�8��O� ��K��9H pIeK�RHHw��Z�3����=\|'���yDh����<}1!y%3�8��:�l�ɛ��Ҙ�V��3��;���8�fk~Ҷ�[CDD@��cj��͸�X���>b����*�<�ЉF��I�H;|.G�l�2�ZNA��]��g|��5l���M}�J��vN�_<>L"{�N��I7�ƛ��x��䩴�2X��Hj�_\̉�@W�����HGEh��3�_1 ��g�ԋ�<09�)e�-�â�=�%��=
�C��6����4*�l�5D0��vo��f�~[K��E��|��%
�	�1��x���A�Sdv�{��5�i<��j��(�Sd��)	f�����*#<�YOJB�$�G���H�Bm��Y:�C�}�V�|�k��oǊ�������q$�w����M<pz�+]��l�z��+��֚����6�9#AA����z��w�^�Z���nYRF�(��p�t]}��
Fc�Y+�Su4m9`|2��֔���XF��￟<�fjgI$�pÒx�O��k��CkFp���%J�PLCZ]��j�jz�$�x��v�F�SX]��m�	���z�A1P6/�d��{�#oi�B�@��w�z���U�4�Q��"����o;\��ĉԈh'�(՚5l��q쪮WW�,^�y&ekv�x���D_ȕe�Q�2�F�0Ǣe'?���V{�z'2�]��J��A5��s�j��z�&���YHө�S��j�$C�;���I�E�1OFs}�F�>�+�A.ͥ�z_#��M+"���v����؈��ԗ,�ӫ>J�Z6Xm?������n��h�<�/����(�B������$�Ӵ�`�S��j�(n�����k�A��'Ah���d��Tt��WK� 2ߧ�������WB )&
���0u �
����4�	Hl(	�=
 �Cek�;n�:�v轨�ƉyR&��^�;�E�B���~f�Q���4�͔���ful�2e�,;N�,��&��vI�#`3Z�d��B�{���Ġ�qi��{'���[��*���!�a?��l.C��Vs���r+�i��ₙ��	���<�\��2�ǕXĪ< �����׀�����[]ǵ�Z�@B��-����F7�-y�yU�Nt:���� �M맍��\�۝�a�1�a�Z��q��s.l�:1�A��&Hlb�*��IJ�֨��y�X��T[���TK-�WFW6�Z��^oiJ��uI�����ng��gOn���~��;�y9�q"`C\_�c�n�������MN�M�8�b�{#[��z�������M9z�K�,Un>ACw����V�3�NZ�#�	u��2�aUd�hނ�zx'V���9�e3X$�����˟����{n��#8���p�N��Y0���&h��-��:�<�Մ�ZՒ�3��3_�R�������˄�؛��TxOՋ�Y7���2����Zh��ၤ��c�PL�$x�ޜ�bX%>h�Ɓc����$L���f�;]�!�y�z�A��nIҧ�L߃�9�>�t�4�><u�
��i���;�%J���~!�p��v��=+���-�7J�"�yٝ�B����u�,�6�4�3���}w&�tP��g$��8u��m5��j�yH��'���8f&с����ϻ�������/.w<u�Co`�β���]��)&f�˒�� A�^�I���H<o�Kz�`�޺{к�5zk�eV���Jg�=��95��k]�gJ;m{oK�$=��iƬ��6gouV>�-(&�� {��.z�:���F{2~3�KQ.�`���I^��ֽ�:���FՎP��Ƕ�`�;n�.�0H<��9�K۠�]�цt��2E��|%�����o�B��j���!�[�딷�ΈYizۚ�h�ڧ�p_�
�����������\i3�;��L�R���ᬷ�����1�1Vh��e��\@���} �ly�!��*�9��[�?���Y��gC:��B�S-F�н���[��|p	��,��u͟tO�_���XUN�ҡ�v�����As�#q��][u����+߲��ΩN�Bc����Q@~�e�o�M�ʼ���Z�����)�74�!����\��=Tsu�1v�шp���Y��#[����5��	�5��-m��K���γP#/�=7MT�EЙ3a����� ��VF7�sŗTg�"?�C*m��?�Vl�Q
�C뇝���=I#��|�%��-q[P׺����G�v�)���{�8h�O Q���=�.�Q�/-xMLrȚ��̞�Jb曢�,��FJ���ӆ��Ls#�ĺ	A[�u��k��ea�V3<VQ�OAW!~4}��e�G(�2H�E:@nt��ONm�4�ȑҽ!{�n9�j��&��K��}�Cm�Je��F��OL4�L�l�t�1"F0�2��Ǭ/��s���\��+��ǥQ<t�MGO�r��4P7����ci�g>3M������ªy@`���*O9���d��6�$�3��n#�&�7���9f�<�{_���pL)<���V�x�� �Y"B{e������1~i�N^�r�BX_D��v_����ڀ~{��.D��}z��>���o���A*S��4�����[��-m�kP�R��BN��k?�Μ��wO�cf!5�? *���
	$�	y�+@D	ev���t^��[��'A���!�YE��B��.�<��a�A�z3}-w��]����U@?$�N!���w'��VZ	�Vk\��7�����x���W�=;;��~��s\y,���7 �Z�I:�}��@���v�"���k=+�d<o.;l1*��e�l}��+�V ��>*�4��m��O�b���-���١g�[�V�����^�g�|�ڸ(��J�)A�K�zt�l���r��=��Y����*�ѓ�^��B��2��(��K���r��5�xݻ��7�L�Hv,��s�SXlOWu"��;~S�b�@61�,��Oˍ�˞B1�g4�����hBe���&n��Yvn�A�CL�7��ؕL�h�Q��]��6X���wd�!���p�D�����;�Ov}"�n	J�o�fVd2Gzͽ�So��o�^�[�H�O�D��n�?!^����w�k�[���a�<�A�&J�;s<��Z�Ok8����I� ��3��>�ϭ��q�`e�'�as��z�u��N�Z�P��>�#��/q�	Ȋ�U�r"d@���I�B<���E��0�S(M4y
�Y*�j���hI��<w|�>����f
 ��.Щ��j� ,��|b�6�����7�\S�U�z�ͩ��x�����1y��_���z��Dl	���Ʃ��O��ĝ}�B�EJ_xr.��A��$[e����}Ӏ��q�p^Wp>����)��������j+4H�GW2A.�>����"�9G���n��XY��J��@�)_��"�z�MҦ����q�����E��,[���u�gB�W�K�\�J���FY��5|)�/ʿ�d>%E�2MV �䁏����8N�Z���M�2ES9���0�uv��"e��(�� �W1�%��+n{���}Wh`TL��X6�#'�k�rl������&G^(@��]S^��v��A�H�O��A�^�hl%��Ik��i��Q�3
m�Bs���B��Ҫ/��"N��bY�x^�m��t����A��Iz�>\P��O��p�boz��I����lp�؁-��e���@��}��C��^�R*%�$��WC�����+�J�Q�MnV�<e{�y1fD��A�QR����7�4-H~�,հT�@�*�H1��m]C�6sΣ�s��
�Ն�s	o%:�4=\Y<�����b���<d����B�_{��솹*�y�֐����x��d+!m!Ly���zd�s�Du>�Q�Ȫ0`���`��	l��_�d�X�ȹd�4n#�XiRθHlx%e�u؜�T{/�ζ���'6î�����ӡ�{���`D��!�f��P�bG��*�MYp�}#��@����Ψ��e����`U�>�o�~��Q��}I[i���w��zD�/��M�a΀�}�����@�𓿍�-�o}�o�Xms��'4Uڂ/7<W�lseÊ{���=<����'�Z0+M��Q+I�Y�GR�}�Љ��݂�A&�]t�]$�"���"9���:2n�
�z{��`��5����:�g�6z�]����zP��7,]�ާ`�}8���3������r�S��fi�p�� ���z������[��(ٚ�3;�2/�v?V��3�T�@h�|�yŢ�����˜�tx��8�)\	UR*�!_�UlbF�[D��g�×1��6-�d�8�n�-.�g&���5Mø��.� �_��j�� '�UZ@H2�x�V���
�y�A�:������4�X�r>�@�}5F#Q��uZ��R ����7�M��ܓo�}���$Dp�WC�Q�k&:�J��ȁ�30}�mr�8����[������
 �&�� ���=FE�J�qz��E�|WkS��A1��<��co���r}yɽ��wt�r�ٷaA�d�����|Z�Q"[܆V����Jž8�A�Ԯ-6�p�*�[!MZ�m�(�.TaÀ�^�w'��x^��2:?V�c}G9s���@�@� ��m-WN](�=)D�RUdp����Pl��6@~)��'�]dD����+⃒N��1Г]f��?�o͉��~�&ҼR#ݡ�;BRm_I���m������j:�-m����|u�Y�U��/��F�DfB���/Ǻ��Kw�0ڀN�^ �f��~C<+,�.���lPO���~f��J4�Y�>�ƶ���O�3��E-��]N�569�D$��S�C�j���*��?8�ig��`U������"�������q�/���b�$�!�G��յ��t[&6��3�ڶ���~���4�-�A$V�q�z���\`���߈�)�K����@kZ�����bYs�g�7�iݸ�O����bىIȫ��VB��ڈ���>$��b��:�yW�����L��W�{���j��|���޵C�t(�X�HXS���H�wN�� ���f��؇�\�	�Xa���;`��]�]g�$������#k�*4���|��1B0��Q��'�d�G���Lߵ	�=��l$&��xPI"Y�.���X_N/vv�\{p>Q3Ue�Zl􅓣&��!��Q�e��K6Z��D��k�����T�36{W���qR������݁%YA��qe�;��������&N���n���7Y�V�$��}���ğd��K
�S������aV���1�7 �y�89��}s�F
��4�*���(�1��/�a�!C��O���qp���X�A����{f}�Jo���Y�q��j�`ӽ���x��g�B�/ˀ&|�	��P!e�q����D���&��H�4bq~Ɩr����;j��I�qu�6�p��Fֹ�L�;=�4���鸝�}��1�4�z���L	B���&���
5w�2��=��fsP@�	���V�>� *�y�֯h����3G��,��ᏺk�S�Z��#��%3��*��W�?���ZP�K�k�o��_�4 	��A�T[�ã="��@���+e`e�$���i/�姵�4i���[�V�[��.��&�p��k�k�A�����#�&a�Fⱙ(�/�0l]�_��Y�G�aF;*G*��?w�w��װ�ʣY�ܤ��3�G`+GѷP��)�N�֎��{�bw5A��c��מ���'���8��^�.�UVY��a		����c%�\u�sB�ؼ9-��^=�״.�up���c�̳=Ϣdflᛩ/m�����O�va�k�0���B!����@�	.����t�e=���U:�,z����pΊ_\�0��Ȓ�]���H�y��+�KP}R���?p�-PD��M���̧���M�wy�u	��wM�8��	:6�".<�ZR϶e�N���\i�_���\�Y.���AJtAξ�'ޔ����j]���]���H��iP6�3�|�u_3:����>���jU2?���P������|Ӿ>��T��S���h�5��3�e_�@oHqbM�
� �>b� �q$��6В�v2i�&�հX��+�+�Y���<*A,U�������>�C�K�|�Ńe�Z��?�epH^��ps��tH��v��3��>| ����ux���W�������5�����Ǫ;ˊQc����ĀUmr�Ј��y)L��e�l��Ke?d�yԻ���tWz�'~�t[h�I*��0>��X�?�pƥG�n��$�ېp��FM,�V� ,<�-�H��[�!h"a1�W����	���3��q��]��M,���ݟ%���y���mId������s5�X���"p���<d�J`�E�s���#�[���i�"==I�ΞU�l;p��֕�{r+���&�]����F�O_כ�����+���Z�A�6>��⚫n(*���@����O*��b�2O\�IV 8H&-��G9��UΆ�R7B�sL(��]R~aB�Jt,C�ʉq��+�| 
GenY���Pd]R�$����u#�-�ќ�]�lR38f�1Krb�A���c��nO�w�������u�=3�f��Z�V!�W��[2��0�$V�rm�� 7��x^"�V���NQ�Ş|�?3X��m�	
RX)�l(�w�
�}rS�,���I���o��O��s�8��*�Zn5�׀���<�J��o)���EY<e�<2��g�	֬�7��˄1~��#�e�W*H�>�(N}���O��k-0 �®R�X��g�ͮ"�B�mC��M�ҧ/�$ݘ2��/_�K�8��eH��-�&*�g��#�_�OVf���mڱ�'>z�?+��gi�mDŇ�W�;��۾�u��G�d@ճ�(XB����]��G\Y�^��|��1��Y쪸{�/�@��,����X���dK���;\S�qi��G|���}����"`�`�s��R�����G�wSa�+�ҽ�ܾ^Mǈ��S�g�o&�L������������a�LN��N-8J�W�����T�Y��@t|&WO����/�c�&fvM&У��gv<�e�k(PF
>���m>%�ȩ��̳��+9����,�A��3?e�D^�W2iq8���l�0le�|���Fa¬OU$q[̦��#��3r�$��T�4dD�΂r��<�Vʫ}������qF��o�?��2���"A{�7�=�h�A��/�F鵡��J����[�_	F�����u�CR��2�|G�2��[+6kN�����m,���R����"�A��Ixg��Y>bAjr=�FH嘕�Q_� _^N��@s��/�WƢ��F�5�t�J9R��?Y"��	��14|IqnL�c�Xx%�[�Y�`������O[:r��;I�	k���f&���SK�����F��������T|	nC |���k��h�q��6j��Hk���2�L�)A����4M2���^5�<��,����'c�K�nϱ(�hc��9Ր��_!F-�?�oW���+�=UO �NS|���Ra[,��ی�z`_pV��e��,j~��3TO���p]?.��(�iE#�^ $AM�x�|#t 9 k���kmO.��t#�y�9
�c�{o����ۭ��@��S{�>tqT!��e�W��Y�	֑��q��ӝqba����t��q�Z���u�ǣy�1@%�Iǯ��%)nJb��GSZ������S�%��J>hi��X��pT�y{��M��Mjn���F�j����/J��l������ߒ7�v���a��~�� >&�ﭪ/� �:�U��!��t�YS�~n��4ݸrP����^QAn�OD�Ź�4�󺀓��L���a� C�+}!*	y�#g����-s���;�<O��R����:w�g. Z���1x�?f�(N���bV�O�b��5s����"~G`��$*
�+х*J�	�C���s�V� �!	�gIw#�Dx����������A!og�P�䑩JN��zز�0e��	�ן��ȇ�8�ox�[�� ���65��/�j��t���7VG��eFOE_6�\���3����V����Y=d\���OâE'$�M��I͏=ֵ�+�K����GA"(lg7=k�t���4�喯O+B��}#I��ˑͤ����Ђ���� RdUw_�%��S������X|ev1l���E|��E�e�OP=��;ø-n�?S^��GĦ8w���[���8�:čϠ디���*l-_w��X̾��kS�$�9��X���t����!f)c�D
��K�j�K+���'���?�G��ؙ�!M��3��IXԭݼ���.Q���&q�?|���	�M�>9�ϭ�����=v@�����\�ŧ��ul�0 ���$/8��[�!�i�эxɓ~��m��u~��� ��~Ak�s�k��g�t<az��ʅp5h��V! skJ}OµH���̀*���������;^�b5�h�����jE$ƂX{\��~(ܺ�qD��x���V��a�J���0����I�y��4�E~%��#��F��[�;��v=$��Y�dY��z�;�wS�L8Yi�{�z�ጒ^�~�pAb�t�)ƞ��m���0;_�#�c���v�:�o���p7��gq�*`�`�\5)&w�a�Mty�sr��H���}��eC3Wom���K��2�z����j� �<��{���G-�|h4��qI�5p�Tn{�oehLd��r�ƮT��a�*ܮ��,��84w��R�է����K!�k��-s8�h!<<ɡ[EY��#��N<�Y!mm�A~%��hR�ё�Y����&hT�f�n�)nPe�Q�=���i<Gc�i����@a��ny�H����M��Q�t<���z�*�h�u�9�g ��G�]O���3�bH�ox��f�/Q���Y�Ed�m#�����/�K����Ԕ>�٩�cL�/��K�����m$N�����5��� O�lAq+G�q����|��4p���)���&w��fJ��S� ���t&Jm��e��.;I�!�#DK2���=�v���tL����9���f�U��(e�?����mՈ/@ڈ[+��Ȏl _��-�,w�0�>x�eN���6�t�6g���Vl}�����d���eg���]C�`���]� .�f�UY��[�œ�̓>uѦ��ҩw�p�f�kot�#D&��I-�9z�N�u�1k���)^l`:���Y"ZNpw;j�3����m�Kݯx%�a&��PR�֛����	@��I��1t	F�)�m�p���В^� �Ɉ:�E��U��Z�R�~��Ba$�#.}�50 ��?&d͗�I�Ւ�c�믘N�&�{Y��M�񒁪����c�B�����qY��_�΢�$�Q��	)�Y�ڂ�e�	ޜԆ�T9�����s3�|����<(S������~����j���Pe�d�+�I�h�{.[v�~Չ?&Ђ,�M���<؃X�$\�t�����@j���ƻ���1ӛ�{)�m��R2�(�4�=Z�/��iv�j�'Mg���ۗ�Ц�#�r.9s+�z.��ؕ;�$.�`h����u���v+ڬ!Vf2`�=I=�Bh�>N�y8�M�����' �/�렑�	�Oc;��9E\�:��P��s����5��Eo�A�,c1��}���l�PC��3O�o,"l&�ޯK�vy��ф�|v��
�9ғ:H��h�TO)uK��DX�s����@���6��q��+V�{��R���!<PsF1�-��-�ql�ɩ���7-���޻ݑMk	��<�	�-/��d_]9.��UZ�<�=dU���H���1}e�d�/(�
L}(^얦�^���QeXYJ�Ң���GT��	����gtq!�MD=�a�Po���!�Θ�ho�i�f�D�<��O�nu*4��x��0�*}�ZO	%�8����=GrQ6D��a՛�p�͌��B�$�����3��v"��$5W)&���EjR"��+�F�
�����-?�'@.O�|O���� ��i���3m����70w�fC���1�7L��&��������!�./����}�����.�ҍ�U?uO~�3 ;qzm\l`&2��G�K''L�z�W:�^hH�Wg���]����(bdp��<�~C/�� Nr���;���z{�"s,���Ȝ�8=&���!�!̮:�A�e�47$7\�I������{Y<�Y�@��4x]-f��/p(f���`�C��.��Р����;�25�PD�)#z�g���<��p����&�Q���k��C�+ ��<�Z�˃���2i����U��w�*�<�hׂ-?4?��J��N���먁��Br��ҍ��~ooF!�z'�5\��XE'yI$6 ��"=�i��`s�ӋN�ewh`�w��k�d�#���t����f��i ���ѭRT#/�'Hb�WD8
2�!���{r���x��;�o�[{�O�@߷���E<��'��|v�<a���'���O�u��V9k[ܼ CL�q�vP\c���~� �<�l��;/�M��Lw^h���[*C�:��l3%�g�Q�83�M*�;�`����b�b���ş��;$]���g�s~����d���O�sK�3���rC�l�V���}��U�w����b�{��#���ۿa�k-��P����b�Ͼ�&57"��%�/n\�,��C&��6��Ppt�w�7���A
��;Sc�w�Kk�ٱ`I�x�I�X�7��u�[sc�?@f��LF��(J�3�i}�%#���hM3��~`������b�pv7�U���N~s�"F[3�8�f��9L|��2���p�xrYlgA��+�!�܃%�U�(��7ok���[H�*�{��+G �o	?�yy��8λWX�E�g�
�c-+�cu���R��%Zb.�5���h�,��ؘ[%:M,����1���h8m����h�^����O����R씪o�(]����0���Y�-����vN+��q�>��[�Au𯁉�-Ů���y�6���}���p>��Ul��Ј���y$]�����#精��yD��R�*eh�#���8�N�T7u敮_ų7�`=��KV*W��־�&8�2�tn��w�v�F~���A9�.�6�0DBOPz�H���ԅ'��n��
3�8�k8�2����
��ֳ�澪7����b�@7�ƫ}0.f#�&�-��
����~�m�N)!AS���}#�ܸB���.�cZ�oQ
�~ދ�������9�������\o�U/$�o\�\'�a^�&�}z��25:Z��<����ދ&P�ZϡX!�@�y,�f��.�\�M>d1�t c&;T��*q3��V<��qG���wf�8�G��:w
a�L�z���*kD�k��E	]��}�=�t�G�y�:�=`�ύ���A�s�KK��� U����U3��D/T���	.���tu1�0 ��a�?�0$��j�i�H{mP�GЄ��.�|��3H�����V:�x�h�0uˊ2?�LV��k�g����g�"R��i��X���G��)ҕ?V����2��b�o�������c7��y��P~�ֿ��8��ۓ�&$^���d��:���+���19�Z�?��Bm���c4����;Ћ4���XK��A�+��*�Ϸ��s�������ԣD�MTLz-G_|B?��ݙ��끔��)b�~d�'���s��%��<r7$5��tʇ�ս��ڈ��usR�qm[sˀ�/ ���(�Zg��#H6�V���B���:80���;�!`��<�胖Ր�Q>��	���)�󇃭�(�.w;Eo'����ԋ�<�����EV7�0�L�,��ȗ��D�oaA�|������������l�3Տ�D��Y}y�@��;tRV5E�Mҍȱrб��G��،�����"-L��`m7�cG��(R�#���znNPWq�,�k-��dyX�$���Ѹ?�O��.k��׺N#*2��	8��}���絃�A��z�B)dY�{�ޱ���-~~D�E'�������-X��U6�l3�Y�3 .�x��K����R�q�{^���Ѧ"g���\)�K��h���ws;[��ʈq��������*�lI���X���a_�F�C	��T�i���h02źlz�C��L�,������� �䝩��XtT�j�qZ���z>_|��rG�ZJ5�Tyزg��Feߊ��{�.5@9��=m�O�#0���p��l�ΜN\�.JC;��u,�T'��G���"4X�o���k�]�����):N�e�Ij81f8�[�k�rׅ����#?����.M^u�yD� �!�7����6ܬ��ӥ7�Mo�O�LtZ�U� �a%8R볐=��498�%�l0%���^��H��#l����M��y���W(����#!���� �tjO�|{B���q���K[c�/=w@�5?㱰^'���s矴�j�B�sg'*���h�[ ��P>�~���UO�1��[�8qV��˄��P�ȣ��ݯX�b�,.��y� �m2��$^A;�G�����-y�4�#v�8�,��*� g��Ĭ�5�N`�1��ʯ� A/}�nH�&�slC�[TؗX�N_Y�q��XZ�/Ѱ�cL�=b	d�^!
pՉM|M�)7��F�!���Us9jJâ�]s�vH��i6�Җ�yAenW�Ο?��zn������W�?:�6�<�'���ߩ��Q%Y/ф�T��Rn7c*H/��o�ݑ������SX�1F���	~VE�9-7�x�cQ�'Z�_�c�����$R3#rŎ$nTj0�g�ʲ�4�(Kۆp$8<��9v̳ޯo1�^�M^�ݲ�AD�2T�k�����ǣ��Le/7�m�a�(�K�:3>�s.���"0~�vb����P�MmR���Q}��H� ���g�e��Hi	��X��cT�c}�6�B{�+j�Y��ɣ�Ϻ��8gJ��E�GM;�6��z�5�ﴅi;�xl�u5�__P�xb[�|ʞ.{���Щ�F�D���E�⟟6�8���u؞�K��R��͋	dzq,��b��
`j:��F����k*Q^��3��q�aR�	�����xh�w�6��e@�_�d*ă:�!T�8��&=�Y���1���0�L�k�!Ѱʂ�Q��0� 
yG��&�w��RM���ĶB+�jU�bS��*��Lb�6��(b�5�z��◛�`��
�����|*�x��p�ݦ��{'��S�W��u,O��d�łv�=���\e���m�$����l�������J�����/?t���85�RW2=(/�e����>C-{�DQ�ƊEbd�p�t,� ��q ��,��ђ���,�&貙)���߱��{��)J16?�	H=�M��տ)Ǵ���T���n���m���tGasz�r��L�y��|z��|=��T��\�4b���C�<��X��o9�l��~�|$GJ_d&yN��;�h[`�~05lCR?ҼvL6X	\��`��"�ѧ9!Z-|�k�rM�!�/��Vo�� ѕ��d�q&4' .K�"��p���?Ƨ�a��"�"_��7�8����o�T�e;�8#d��xAOW��U1ȇ��c����=�P���3�+孰� �@�(�rc���(^ �f�d1���n�;��:1��6A,�����&?]:��;5��mΊDX*\�ԁ7�Jwd�=�$;4ȝ��V�t�K�.�~�9�*�9ͯ9} a�3S@��	!�,x��Ug��>����($��̓��u;��!\��UZ�(h����aD�|G�Q�V���j=�r�*ۆ�uC�>����k5V[�~W�d!Wp���iI}#�J� ��efiGv�!��B�ẇ?�J1n��F�㌤�[�s\�,G}��K���?�EK)��%-����PO�Q����9�'p��_e��e'�v��v���[����8�*��2f�%3Er�J~""o�|1�.�1������T�|�#��k3�x��+����0RY�1���|\�W��6�N��	*�\�S՘!p{q��vd���.&EZߌ�����-�J���%d_�m�m�������V鏸�~����fڿ�+�x���%׸5�ƽm���Ǘ��&XFoeVb��F����%"��]{�S�QN��z�v�9�`&9|߼>���(���Φ�f'���v���u�����FP4��Q��>�@�B��U���=��w��쇎��"�O_�HQo1�k��S�$�oq~�Y0��'�^�q��xء����K}�B��(!;0y��-W^���IM}�!��KkV*���������cfԻk}%����t�4�ɉAl�����i���`���(�������I�i����F흺���|*�����9i+#"u�0g>YZ�j�k>Ex����Y�~ߙ�+�I̧�N4��O��ߏtKі�z�_a�"�)89�T��!P˄}�KI��x�qI�;b4�=�=���X��YA$[���k*}�C :JD^U����ĶC��ֆ��
T�km�l= �j�
j�����e��-��]aE�VgC��	�<Qi`��	M�D�-���=�G��)fUҤ�V�^����n�#wy*Y�6����ͻ>�D�� 
�ρ��A:)ED��i	� T�D^�D,^���fܯjP��Ի���r�M�Yg��"��o���ziy�ݮ��uDJ��(�b9\@}��L� r92L��@��Ϥ#���o'|K���F��֑�\�C�
p�򼇣�[�E��CƁ<����}�A����Z�����e
�Cd U�;r��#�/�W�,"�kV�����L�W�����N1�z��6X�"}X�����N$F�P��"-��J���G�ۏ��Ih������K:_�J5m�H$����y�y�����0~��B_�?PL5)�����(x�|�����x��*���:�'_�v��Y�&�TM�84�o�E��ַ�>�}yvSN8DjDb�ۚ\V����RU�����f2���1 �qd��<���"���ܟphT�f��jN�C'�6{%8v�?�G�����'�u5���Y8,N�=��y�@����"b��z�`l�1��%�V��*H�P*���J���m����KO1C%�y7���m�S�Q)J���X@�l{��WI���#3���P�1�e�
n�l���䶚�cn�J�]ۼ�H�4�ND*p��K�e<���]*O�����@0�Ͷ���$��u�3�
S�'�{O��R<o���M�AC��h>'����i1����	�N��%�vz�x����.:(l��N��<�$p$��x�����q�"��ci�g_���L�*�W$ٛ��V�i�%��������+"�F�ި�w���0-��"�#\@<0����f��t��
�PA�p���+%�qmx�<��Iy��a>s�/���q���ĵ���h����7�?hTP��"�t=_5�+�+h �n�s|���)^P�+�A�s��D�f���F7J}1��K�I=�9�TӈVU��NM��7N�Q�ܦ�7������(�A���1g�������ݭ�o4�s���j�D����>�k=4���`��no�R\�g��|G5���J���EL��+⭉V]9{X:P�	��n���t@^P-��Ux$6;�$��3��t�I�	ߩ6��I^w�G����x@{"h��@i�~E�:�S9���L��]��4:B;m5��q��I
����'���I��a	|A����-y����p9�h�DP������G�oG��%��]c�E���Mmmٯsȕ7^����̔U}�T���)�C���
۾���X7/�Anq-X�������R�IP�`�"��_���a��;낉l�rk�UYߊ�e���6��:���:��	��_���w�R�;j��j$ ��י�P��l���~�A���9ha��r�$6w�zh�H�r(��zr�
#�����*r9�T�]~�b����q��`u?�d�|�Ň��J�M呏 ��x�v�CW��#|p+LH6�d��� .nK$��m2�N�Ed�fXrz�ow
K��ސ�8��g�����<u��;��d�Q�*��c|˪o/tVIP,q��m�}�*�Q�5@���=���k��z�(�V��;�Y�<��J�.�K�5EO���ȓh0a��CWIHz��m�3>mk��Ә%5Ll�*	Ԩ dۀ?!>߲��.C�療Lf�J�
�R��V�{c�Ҽ:A��O� �0X������v��f��,�"!�_����� �n�)P���?%�� K��S�i�o���{��Ϯ�?߫ ���
hj>�q�����K�s�oN��~s��Hq�*=[M�J��	gM������@2^�e��<O��^�Y�n�k�Rr������LQ�ވ�?^��:�P�nO�(�ۣ$f*x�xL����}Ѥ�,�=
�s	o���<-�S�Fx�-��[�4��F�P�pN�	���Tv�\�þ^	�f�h�y��EV!<������ �C%;"9���>?L� +�n�{�|�o����e��W�>�{�E������ư�Q8ޕnnNXO�#WakQ;A�hV���>Q�I��o1��(f&����ݯձ������;��=�D{ �լW���׻ X�ҐSՕ�_pU�S�g�>��'\�:�2$�V����h~?iI�^�q�u�ä���f�uK�Cw�����U$�8�(��>��	���7l~zh������Q�qÊ9�%֨>;m�ߝH��u��f��JY�Q��
�0�\�F_��ZM!^��@��}��Eg�J�ҹ<�H�[y��ǳ����i���6�BZ���'��[q�^�N/���58��a������9�%Җ�b���#*��\�1wW�g�ɣԊ�~��a��:z;�(:jk�dsG�]}������ !�>�t� ��
[b�a-��mW��D�����E�M� �{����swN#�_H)R]�F���!ٕ�� �M�}Ou77���~�A�IH�(��!�#��}x_�n_�N2��c�,-!UYR�Z%V�y=w1rꏫY�n�<��o\����-ۇ�J>Y*o%�Ag��Ӻ���:+Dyfc�.O�
��\p��y�y&iX��.��m��Ψ`��<��\���B��/fL��ԗ���kE���{�}F��C��:[��f�3�C�f����옶�,�F	����Po&�!�U��M�y�'Td&��D4��@�7����c�bnAo�]a�Һ�U���e<b�Ƒ6�$��/������i��f�Y�'�E	�P�~Dщ���^X7
׎O�=�8�wݜ�� �_�q^�J>e�pl_;'��qq��4��XLO\�(%�%0��I���BD˘\��g�Yb8��(���(��e�=��1Gꍝf$<@�h��!��)8������E��ʡ��jy�&���,M %P�mNJ��o;��_免?ٝ`m�5��7���b+AM�s�c�J+i��j��)�8_]ܟ�5����@���/M�O���/����� s�œQmpz㓞%��I꟨��?N`)c)��1&�K鄙������8�4�)��ڇ�Y����j��v�=�'�A�Za�>��������n�c�>4�I5,f�ׂT@O9����ۭ<�����	�1
�WY��7r�]�>�M��v5"�B�K'	�L�bo�H����{�,����k�|(ׂ`�!��٪��x����u��:����/e�>����R�^��
e���|�֎��|˱���f�sA�;�x�Ԣ���E�>͉f�-`��� ^/�r�:"����yrk_g��d݅����Ú��OS�{�E���`�$�^�a��0Q� z��<�� {$�~?��q�����I�I�fi�GXi�&�r���7����Xюfhk||���?AV!R.[t��L$��/�;��n3߰�EH*~4ۃs$i֛�56VEfe�Z���/�t �P+���� �V`�ۋ�$�Ŏ��=k�!��N�"M6��L�/+���1kYkhiS��ΰ�p�nY&���s�H���1�J?@M/�Ynf�Ez��7�`Rb�EX��Q�Z�O#9+Ye��SH]v���WӗF ɭB_M��T��yv�EJ���W����*"���^̿4��� q�~N��/��Ԇ��W\g���Nz��G}
���ഉQ!-�h���NK������ٯ_��Pl�D�a�?���6zw��j}� Y�V�yI��e�3�D��L��AT�����vRi��RӪ�l��w�I-v��8�H3R0_���R�lߗ�8�&����;�D���#�5(,��&���Wŷ���H�@|!�׬wCa>L��ɬ��ƀ�Ak���sG�*u~��T08�1ۮ#����T���c�v����;Lhl0�)v�`��}.3�[]D���HQ�D�)� �N�~/p��rF�B>�?H�J���"���|d�՛��N
y$��76)�Ql��\�Efʳ���Ҭs�Jx��-���^L��N�%���p���?���\6�RE#'�ۉ{=u���&_g��q.��)7kk[vL��8a>++������ު;�8���-'��[����w�_�:��K�Q{621����y����f��A�)�2���~ܛ�?$���"ï�����)��ک�0����pyM�d)�jq�{R�%R1˗�(R�$"�~�I�p�Ւ�P}�I��)[� �����I��|3$�Ykw}u��
$�ŷh��|�����[W��ϩ�I�I� �ꉲ��rH�ז�:O�v��´Qެ]�,��E8;��Fb�ϔ�}CT)'�P���2>s��͡6&�nøV=�ep4䴻��R\;�J�Q�%ZV���_�^p
�aK��
{&P�p7���g���r��,��7G��N��������֥-ep G��w�D&fǔ���<7ѐ3!޲6g�Wg��,�	4����a����f�o����B�=�|_|E���������Z�ց7��� �`=��C�,��3=��q��{z��nLY3P�Ӻ���RK3�8�P嬙�'��/R��.���҃s+�Jm�� \��^���{���"/�O]�����Q�By00����Ƥ�ɞ��/q�L�\�+�>���1{C����??b��&xsx7�ZiD�:�J��޹M�v�e��L�|��G��?JE~qÇ���7e�jS�ȟ-�'s ��A��&\��17�& VMZ�D���P�a������RW^Y����>T��I[GG���/o��;�եC�\i/���K��)_�>�m��T�\?:q��8����QW����KD��U��~y;�|���ψ�w4�8{��3w/��˫	��RT�<c�d�Γ�G���6�Χ�f;m|�4�]o²���E}�����P+�&�1���5?����߮52��!�3�JWo�K]�]]��#>�r�p�)0��`޽]��+\``���ϴ�|}g��� ��\��4��fC�vD���~C)��J�(��zpa/�z�Ķ�f%��ؘ�gĽ�@q�]K��h�ňL0�V�\�e@C�LlV�~_�ɟ��=?���d�I�����0}��r��p#O`,�Ĵv�@P(��LD��k���]��T���PJ�p�i�f�d��r�*���0���͡��,43��j�7�}%���(f�2�B���f��Xޡ#�e�ۨc�,"�����A�j��s�*��i�;�L��j�A/�_�`�5x܄Z�.(���+>�v�ռy������{�Q�O�X���K�
7q~���bE]z���&�jV����]Wo��Q<�8�͖��g�e�HWΈ�1��3b�{ţ���g`�9q}�ݻ�/봎aY����tL�������L,ݹ�ţb3{��N@,�7�uB���H㛴f����=\)��B)k� �]6�����F�脯��1Q�;V餑C�*�aG���CϪDa�Ϳxt�����k���6�w� �AЮ��o����q��M���]򁼧���ZOQai��/�x�˽H5�F�"�a�h^�=ƼIg(�)���N�|�Ia�o�{�%�a��%��{�w�����`)_K�����iW⚠o����GKD�?�ݪŃ�vH����t�^��T��%��c@�}����=�pOdw��j��>��?g������B �X!�J-���FB_W����W:>���p�y�+w�S�ͧ.v�QT�B��":���`zNsz(Ϫǲ~�p*��.��U=F9(���9�=���E�;��.�?6ҿBH^^j�"n*�i_hg�q`Owk��S����V���a�8�'[��?��������_ev��3����].��Y2@�����+Uڮ
lb�!���E�<�?l�4��żf���s���gO�)�H&�p����\���Ϝv�W'�>�~S�wru�Y�.���h��cB� ��"QA��k��J��i
�I��'�Ԕ�7)�W1F�N������yP��@��hC^|�J�
fB8�A�Ѱ���X籏�?xsQD����Q�u�	��"9�߹�Қ����̉1s� ��U�!�~�"�r� qET��틮��%���U,�tJ��;/O�XCd�C�OZ~�;�@���E�0tM�tc2��g�X��s�f�1��ja�Je��h4'��|�Ѻ)�kߧK�C��_9 ׁ�@����յݳ�M��֜k�y��<���6��-�eΏju�~t���_�4�N�3y!�<���D��>}l�?2�1E.>q��I�/ �y\9�g_���~W�D&�_�7����&�\!n�����q��Ѝ�>����&f����C�ݴ�Xe��w��7n�^<ko���B$i7�O���;3e�s�0j^�D(э���mx��ܾWn/�F6riig_����-��q� ��_j��b����/�"��p��/����n�H[��� T��ث}\��:���ڃ����ԅ{G�L2O���{ѷ�)ik�{�����v�yu;l���6�iz"%?�<���х���~iK69���!c�E[B��O����Y�Yl!�X�1}��ш
�H�{ք��X��O_>,ED�h��`�~ehm��++����C�b"C��0�c���������S�>�%*�V/�^NpD#}���Ԍ9a=���[�}g���|8��U[��e�8���Y\+�Y���gSAa? f�u��U�rr�U���ݎ�|y݃�V5H6��(*�
�'�ЋϺ�����c��2�|8t�$ �'����X�D=�&��M�"��f��IY
1_�l���p������^t�3s92�,��'h��Z{޳�X8��h������y����R�o+�	Q��%ʟuuh$=F���xv��|�ך�d�Nzp/���l����D���]���y���E. ������t3M�d��R��É6�x� ˗�����g�����SjL�v�����U1�(�[V��wCi��**�m:s�)��U�����/d G��|�d F����]�b�~_F�P����~�T��.=x=E���8��{B�임
0<_���u���g7��=�҄S m�ڤ��&
�W�ד����e�9�N9�v�7>�I=j�N�+
��wS�Wbp%���	+�=b�%.��&�q��c�b[����j��U���;��m�������#B8�&~�t��]��)�d:�u��~�&��t`p�M�A��Y[l�`�se��[���6p��-z^r�_�O@3�h�2���BT��F�������f2��M�*��[cpAԠ�n$�V@�q�U�AU���Ntbٓ�]j8����@�2�4��3ɢ��'�~ڀT@(8B�V��
2lc�X�Z����@޴̹�O�=R�U1<����Ä���a��X�]��������+�|j[���P� ,����R}��A4U��SF�l�\�O�_�K=�Qࡑ�;�R>� �n����7�w��gE��VQd���L��"�~����MYbI���=���Sf�>����)�̕�)e�F���\5��C!T�w�F����?X��r��mF`�qD��T(�1h��}��������z���}���p��g�	uú��~B�|Б���([�!�t�1Z�����~�G��Q<�+gO'h�9>�#&bW-mP�nC+�e��S�*�Uu���l.!�j��U�G1��Л�f��8	W�O��e��F��!�d��e�˿?�x���@]�\x���4��c��q)-����H�H��E���	�}�����@�\�E��wg�*d,��WU�Ĭ(�}|
�eИ]c�c�56�v[�U���pRt��E��ĥ��լV�Z?��_���gO*��&)w��}�#�((�]sk���!����n_�^H���w#��~�>K��W�i��u��7hk�0sCx�}����x�Sy�F��hlO %)`����މ�
�g�� ��:�Pݚ������Vc���~HI1���	Q������&���Uȟ�W7�8�)kKt�N$V��k�����׎$�U(�O�4�hh$k�Ta�6�i�d�nL}��<�ީؽ�1D���+>ͭsO�C�Z8om3Ѽ�I���\���h������w(|qu�뿀`�7J�(�}���\�{��Y�G��1I� �Ż�zLo�*+��(�%�y�0QJ;�f�� p����0���y�H �� F&�����qϾ?�R��oA`fK@�){��È�E`6��pE���'��FI�[�c]���w�� �L�\�Y��	�9�{�_�YYe��	H�*���}R�<<H5�(���t�"��L�p��t��H(���f�d��J��=F�rD��{��2�����r)���P�,H��x��e�NĪ��2 W�5/K.ycf��wD�Ylww7O+�ֻky�!��Ii|��x����f�,�l�C��݊���K��6o���:Gl �SU��l��g��?𦿻�ew_�?����{�r�W���.S��~���Z~���	��Mvc��}��n�U湮L� ���V,�m���B�O�qP�$��?\�f��/�9��܁%�����"�5#��Y��hH���i���;R(��b����m��$�v�]@-�m8�M���z�O�E�4�l�0 �ʢܗ�y����Y�z�^bH�-�o�8wA��޳A��~���'�T�x�%���c�s%�-JSA��������Ӛb+�g�Vm\�3�9��ã]`?���S��%O|c�ȥ�T�����3��zU@��N�L��ie� �+@T��}�@�h�ݲ�fU{JpN��
��v�{�PgI�7���YmRpD���cѝ�`+M�Ӎ���!���t�K�G̟�������+1x���LY2o�����7T��S��xZ%�m|�G&c��F�,g����wG��9Xp?���%s���1~C��܍O�V���iRQC�X�%Ξ��Z��;&1J��u��"n{�M��j�-,���(I�	�4��kTy9ˎ���m�q���i3�뀥V^*����4�����3����K��>�hGPv����1@w���i�.D���i2��`���K︎�陼��A῎_�B�[�-19���0��W�3罎H��t+�5c�0&��E*Gۙ�	��g���B`��(��������0��f_���oljfY��-S ��?�9FI���J�
Zl.�W�x:&-���7�Ar2��(5�xP��2��+̳Ao(M�"(s%"j�tͭ.h�.���l
=����
ҮN�p���䞌��h>�K�K,<��v�Af�^p�"�M?Ze�,CS���F"�u-�hW>=��fj�У�hЛ{
�)9�uGy~�q=s%��W��fA��35��d��7���I+���RQ�Ng�b�����:�X^n�h��/����w����r�:ҩ��[�+ݒr���|�8߽ۻ&d�/��	�<������a�"F��� ���m���_r5��䒢�0�����-�$Hw��u��ݐ��k��e�o~�%�*�8}����vܤ�˃�I{�U������F�~���V���J��ƻ ��������zI'Å��%�����Ӊز�A{��"���8�ܠ ���������osCmJx/%�������<wJ\���-ׄQ�_��"]��"os�){z{G��:����������H�Y�T+q}h!L�,���I3ʎ���S;٨�+�� ^7��(�(C��_0�@��<�CL�aBr�5;EY��E;�Vp� �,���- {�9�A�߾|�G��9�C�j���C<�+���ϙ��(��w'���3�Di��~��`��m�D�%�ʢE���x�u<4{��+{�1"��M�Z��W�Y��co�{�d@Cw9x3G���1�Y��H���!�ω�a޸��^47eS���G��?�߄@Ǖ}	�M=[�c2�'�[b���Ԋ�B�b\���yQ��	e�,"{)�p�
�_�	�� Z���?ĭ��䛮��!���3�|��`����qb{��qq��$(��Ă��j�T;��;g!>�^���h��'�Z# �(g+!�5+7`Ӭ(N�g���,��q�XX�	�x1	!�)ly��s%���	��8涶s�h��j���9\�|��Z藪q���ШP����4	2�R�u:�#Lo� �~e������a%����ˏ��۩G4I��3P�ɀ=�m��Z'������1���� N#>݉�t�bM�|�4]����Gx\�h5T/��UG7KS#�>�4+�gW��o��Ҕ��(����9�<g��9$L�m�5u�q�aM���k��<�,Ȩ�/�(�o}&dK�"��+-٥�:���G�#�p��N�dj��DV܀�ؿv{�Zd��͉,I'��o�8�6K�A���Xx���EMmQ���?��Gw��Sp�Ϻ�������]��R�4��j'�����2�	m�T�қ3��(b���a�Ɏl
k���Q��G6fK�Իa0���t8Lt��8W0��|V�ĳ�a�WE�`	���1C��'����7+��l�<�F���RZu1��n�q}��_qV�è��#p�;��3%�����q	���8s�R\^z�"�	�0u���X�3:,Q�f�.3LQ=�/�n����2������k=c�Q����P;x�3!�j2Q���H ���b3a���i���&�.����V?z��+Oѹ{7>/�k7�4\E���U����)�+c�0��A��a��d<���6J�������7lؖ7��&��B��+�Z�nv�ˣ�Ҹ.(*�����[V�^?O7�qg�?�B�ي�)���ԑ��eլ=���{Eg?���j��4=���p����;[�p@e�v5ˈ�#�,���V�W�Јc�3�(�p�_����sk��ҷ�d�I�kW��D���E)�?��x�R��<�@ R�[���WN��(M��iځ]k�g9BX֐�[���:�*5uD�7*H�%��z�%�N���Y>�獋�1dW<b%տ�)�U��w�_���[[M<��.K�;���p*�V�/Ӻz'ь�ԩ�1'��e.\��-�|�?�Ҧ��;n�$/U�1��h94�v	N�C��?>�EB�g��(��C��c2F���Y��
*b.�)�>�'���M*�Y�.���,T��LN�'s����#M�ِKE��O�m�s��F�F�&�H�6���S-��[b=ȊO��oƾҁ����ß�g�F���/n]=Pm .�<u:E�hm�?CԼ5�S��;p�v)6����Vo�p���h��;Ӳ�i��]���ws�V6��ҙ�*m��]�
#1J��`-��E ����R����N������&�%�K���kP�XU��oGa�p��U��FҎM�$���;�%��t��p��ǽe�����V��˂Q����kjM���{e�:���H`quR�S㨝�Ҝ�6� $��!��p�Y�J��k�a��k��kr�4G�G/������QN���Ҡ)�y���Ib���E��֘ӳ��T\�=r�8��:F8ߧ�g��$wdaQi��~�T�
�DI��H#�l�A�M���!!m��(t[�T�*ѻ[6�ww�yگ4x�_
WĀ$=����&�����
�	�zW��n������Rz��9\ϳ�����G�`�H�t�}y�Y�\'��|��b�#��mI��y1�O���f�� X� �jY��4���(��Yc�eg�wh�M�o�>"x i���Y���m/�۽�Ѽ�S�����A"W�<�ݕ ��{8Z��7�XS�0\߂�Vo�3��C���^A9�6���3c7�s��>"�M5':Z�^�M?��?�6$2^K��vh�%Q�&[~S�pߏXN�����>ᖌ;:c̋��)r����j.4j�]�P��q�37c2�}���]��Ó���T�B�м*jw��C�8��������� {k�eN���/����*6U��w'��/$���AK��e�wY1E��� ��i<�N��Y��D�=(�S�b��Z����l�;�ol��q���nx�����s�++|�)�7�}�VELNu����!>����OJp�(64��&�+�P.��q��8���F��i_�F8���s�<��j�tq���Q�0��Ɛ�yz󼻪p>����n�԰k&Ѝ%�`�f��~�Y���}���HZ��w2Dۙ�e�7���Ug%]ÒǍ���M�:0���K�^7��d�^@ݵ��m���&dO�4�G:a�q�򧝠g�(����P3��)�oA?��]��f�(7�u����W���]���U4��v�H�X�8S�aG�P_,��Qf�x�y�W�Ni�O8�E�)l�䕓&�7{��>Hp��ѩ�KeM�ě���D���}p�Ą�Q���n�s�Ǹ�>W`��|^	>�}�̉��{YQu��y��N:�ެ.Nu��n�BLzG��[����l(�E�����X8S��b�
+��А�d9VF((�=!��/o���?K���s��N��\���9�*yTЮ��[��bX��E;��vd,y=����,��>XJS
:(\b���@��.0@�3�aM8�Z[�KhѬ��Q�d���� B�ɓ.�ޣ�*ɚΨ�(lr<(�|�J�/�}�U�ݨ�K�q��V�%�%�!�8��p��C3�Cԡ�����`�V����S�)<��&��;fBͤ �0���Jp'LU�\Oy��8�@MCm�uϜ�QWĝ��L����=t]����
N�Կ'm����'ꎿR�-�l���`A�R�M¿��C��F�	��21���)���r|3�`�Z2g�U����s�<Xõ5B��895��	1���yxԏC�����o)Qs��vUƿ�R��<���+��>N�Ì��(9�f�S�,���'0�O� �F��i<�/�Χ�Dz؁�˸�؋+j�W(᳛F{��Kk�߮���Ư�QVsBTh���^۶�jY��lq�������,Zi�+d�eb�,M�O�{J�yn�K%¤_�-Կ�Wh���u�����4�4����`hx���~Hz��TB<���Mx�!���e�aZ��R�$[�O;�d�)#�_uPc���ۏ3�)]}�}��^��㎐����s�D�f�p&a��t=R���Y�(4�&�4n�� ",��&�]V߳ob(�l��.n��򩭁NVѻ�^�}�UjW�u���-�
Dj�CV�S���h���w�2���ߘ���u�Z���D͒M�tQLĨ ��:i��:w���0�@8���ť#Ϗ�7/���q�Zy�W�ˋ;�g?�1 ���!$~�`��f�D�R_iF@�{�c�Ĥ��d���Ƶ�J`�	�o�m�U�T>5�PD�WGF��V�VZ-�֐R�$'NS�&�R��-�$]���S�E�e�]҄���z�VI�U���5#��⳱Zd4�k%y�l��f8���Z!���AeAƶ~�(�Eɦ<���WY�w7i���/"=�f)'GC1���N.�1�	<�"�I��ф�蚘��5	=)܌h��"�}`����m�N7�_�t�v�ǆ���@Ji{�|��E?\�B<[�B�b��7��Ȕr���98�l��Q���9ׁ���'��[����#4}����Ǭ:r�$�!�א��S9;�D�<�SȚ|�GR�ㆾ�)�s2�>Be`d���/�Dq��F�Q�R�@��΂n�?	 qYi$�����K=���>6�v�U�]�x�X��I?T��^�އ\^[�>et�_���n�����}��x2s%�J�4@T�5\�4�dـ!��� �In_��
!AY����r�F����g��eE����ڡEN��9�{�q=y����S7[�%��&��{�N5�@��-�X���G%��ݿ�&0'/-F{x6J0�s�CLBx��!ۿ�dגN� ��IG�#��G�ar9I�%L��(���΢A��+P"���{՚߳M�� �N����xr�\�m��[RGW���a��g�]�9��5����Q`~!�O� yE�Cֹx�]zGж =�!��v�L���e]*2��kac'�C��o�Bq�t�IKu���A��g�A��8���i��JLfs>w���c�@��j�L��4��$����3��T1���Y��ـ�؃�JԌ�s$��T��pZir��H_X��(���|���ĖZׅ�Pl��M��*�hə��_�h� ϳ�9��ծ��S�Y��HOW�C ��0N0��ҦN�� �E
.g��R#�����������K9"�2bNF���.~6��nb+��#� ,�k�.yަN������a/�o�a4	���؟��׸8��8�?��^�2zN����ِ[Ƈt�j�Q�$P��*)>;9�C�T��woWM��M�u�Y87��q� �T��@+`�Zv�fc�=h�-�1��hH����ʇ[ƀV���N�P�,�xu�@h"�>�h���U����CZ�S9\� � M���^�����Jm qsM��Rw��0������_w�X��];�짦�z(�eA�yG�p����C��� �KLǢ���_�m_�œ=����'�[s�<V�E	1��� Amɸn\���\'�;�Q�Ȍ	,#�2�w�e�f�Џ��űez@��G�wʮ��Oت����回!c����� �[�Y���tAW��Ni)�%�P��T9��9O�k>$XA3hzz$�O�э�i��`;u"t�?�P�D~YEą9���4P+��h�/a$.C�������`����fV��%( ��M[B�(�M�
N�,	�T����|�A{hݯ�5��'�I�<  �{Ί��o �C�F��t�������8�&��No��;'ٰD�eB�m�У��E̊X����`o|~�Q�D&ra�B���[�&�5T�憑I�;�E�yR�V=9��� �Y�3ܧ�������/�z����Ywm�r���HT����&h���ގ�ϴu
~�i'߱ 0U|G������O�D�;��$}�����Zp"��D[Ʒx�y��Ctx�eL.^�8�����
��&�!���m��:����3u]�	�Ո�}+��b_>q'	�>���w��3�$*Cd���X�z�bB�N�cA]�֠"8{��v�Q�hp���;r	#6��[@�%� i31UXҚ�c�Q�7A��H{�ӌX�BXѧ��>ml�����X&ȱG�|]a����ɫ��bg�` $/��}�M�P:�%��%���ٵL�Ԟ���]ş����}}������7���È��ؖ�%�a�S�x
���j=����I�V�`�4��4gu�D��<��?n�FRk�0U�����]���(YZ�X�0��é!��.L*M�����_�`MeB�)"���6�=�$���rjF�fP�X&�����w`WF;�Q�"��=���W�[{���j�S�G�P�wfl��7�9�5W\��e����`�k��A��7� ]�N�g�m<��)z�
�@5�����T�U*�YVr�� ��\��̗>��<gU��E�.6h�,2�����̴y��FT������-��'k�D�����B����}�I��&ӄ\��A�7�1]���Os�p��V���q�ڕ�@ҏ�"c#a�%b�W�H�]��#��֫��Wrdv�&H!l9�Կ�SW(�;ҷs\�F�:m�bc�B�?`��k�h�]�[�[�p�ĳ'2CRV�y�z�1��؜0��Q�=qU���'����'�!�=�~W���ҙ�5*�}
������!ޞI���|�bʻ^��휚!;�D0e>k�����:��wĪIϰ;6�(����q�ǩ��nk�� ��u ���e���I�ܷ�EP=�|��G��i!������=
�D����/zZzZ4~9+`��>� T��;�9�.�e��h�nF��E���ʌV���'�K
���@�娨d�GJ���y�Z={�B
���d����r� jd�+�a��lh��Q�-�L�����ЃYd�� �ϩ�U�.ה�j��ty�1�<H���^Ji� c�[=��FLՙw���F}54��ݎ�Pʕ�7b��6V��Fu�O9�vy#�+�(���
�\hG�ڨke@��/d�mY�G4* ���PĤ�~���X�h\�
��zw>i��U����L��d8<c9>9C"6A z�V����I���g6�Gq*�o���N��񝣦r�Σ����L�7fc��V5gd׳9�j>���{�`2���v������z���r�{:���Q���2�
��+��N�D���z�>=ȷ��ਵ�xf.7_�1���3j���{�Fm��7���+T�%՝����~�WU0ww�n�4ZY���X^.�w�J�-�	~���}����=\TV�.�o���H?+61(@�]ǖZ�~�/x�$�8�����k�6s�J����}h̆p��L4�_��ۨ�[��{ ��
ֻ�oh+>!��¼�kEx�w/��q
���6k�U���~lA?|�@7�O\�ȧ�� u�7���t4�w�DR"xm+RuB����C*H�)*�>t���x��zݤ��f`8�!À݇���JL�Y�K/*DJ۪�I��05�Bcذ� ���Yio��5��Y74>E���_&���s��'�����dܦ�h-�F,������ᨨ�7+�a�hL*!R9�X�)-~w"XOHq\�嬖�~�4��|�����ԭFK��I�๒Ɔ-q�bu����KM8|7�����'�?��MMP�������z�R56�0�.��������*Xή���3)[���2i��Ü�>�`��"zzgo�8��U�@���[	�v���O�i�������� γ�q�\�f�^|U=5U���vM$����*�V�M�j0�LO^�:=8N���v"��vivL�J5js��G�7o���|ꐡ��h�?7&��f���/��lS0!�X��|D�n7���}c]b�k�v��7Rn��Gk��N���4� �Oɳ�j�@�j(�E���|�]1��)�&L��?�0mk+ky��m;.�0W�q�>�CRo����� &� Opm �{��鉱��U���f�	<N�%r͡�Eٛ3��[�Nüa��U��׽�����CiRC�ܾ0�!/BP4"��	��1��q?�`��� <�����lW�K�!�I��6r4PIi�fœ�?�a��2$A��
������<W��M��!*���ZG�S�**HĽ�@`�j�6�oP6 �3:Y�?�q�!f��]?V�o��{����P�#}L%ޗ;`a|�$��#�M�+�:h}M(凌Ȩ�L;���J�/���Q��q�.��Kg����r:���Z�+0�&�XXZzWk��yBw��#����o��6���@mE?ݥ�/�b�҇��R�{��p�R�y∐��&!#Ø���b�B��[�F��/炡�J�q��%���l�U����Ԝ�F@:�r��'Ϻ�k1���[� F�
f!���B6�ؾ-g����C5!��W�@SA�s	��^򺉫�~���b ��b�Ŧ�m��QP�t+P
<�LB5�q`)�i��X=�|��*����PsJ2�w>z�!��ͦ���@���|ZR;�iԍ���� ֯�B#L��'C��"��C�a�n�R�k$��b�N����;��Pg��gl��;䃶^�G���D�� �節�U/��z�O���V\ߘ@^T��'.=̿�H��m���m���YB`H���4��6m
�%$(<%�F 0�D�y�c��a���ѫ޾s��h��#�c#O����~�$�Z�r�ֆu�.ʞU�%f��2��A�!Ή��Fn�����o�<����gw������$Q��Y0j����&:��^[r7�Id4�� ������d�Tߛ�?ޘ�w�P��?z/��B��|�/����Ō���x ��"�y�����(�'cBՀ7��0Ҙ8L�U2�a����M����A/4ԡu�꿄����lR���+�jy�U=(86ٌF&iա�i�	%������~b�>���1�a��o��h �K�AK.],�	�8���˟�!���]�ղ��*9:K�v�[��6�X-)�7~��6`�'�/7�n��M|��,ٚ�/)��0ɀ"d)�Sg}B�rR��m%�� ��`�lX.kua�:��Y�_�o�2S#|��2Km6���Q5qT�eg|_K�5C�#�C^f�۶�nr�փ��V��m�1̳���X��>V���ƴ!;�"��W9��l"6�$�f���wrJ�^M��.�Ò��WloT<Y���&�5G����=��>e��T�UR�+������Xd.GuIJ�ya��U��/	C����m��%�]���S��(��l�3�1@ �?]�8�=��*.I���،��=Fǡ���Y��!d��g<�d6��,���R��LI���g��ז:(�#;�P-z*�4=���i��Ѹ�c綷M�eԫ;�U�R�$�!��#�1뎁�Ή���z�13�D�J)�����q/c��V�C}���2���i��{�{9�)m�X�����ny�����!��Nk!v �JQy*L{����/	$l*< NC�R��kavTP��=FwJ�`Nc���QEh9�:�iI�;P�I'�f��f�*�`�)���Rli���������gU��}��W�,�g� �4��
���4f 4��ƕ�I$ܕ����
E���l�"�~p
j�D4:8B�Ap+��l���a�)F��q�]32�N�<��
��)���\�:/n��+Y�����4�����=w�P"���@-���:�?
�0�7۪�_����gnH�E#��#e������o��-h	n8��%n�`��Ԭ���K���2�/��j�])#IJ���/:����Ǝ�!(<$\j����(t�_��D�}�����R��U��R�nL��6��qrC5���k�� �qǓ�b��v嚎����"f��Z�حT��_�'�;g��g��˸�7�؄ݡ������1��CRԇ���6a`����%��� ްq���5P̮�+o�-����ȕ�~�2�_I��٨�������l�3�p���#ܦ�j)B{eA�MX���Q���'Rd�T�!�B4K/�Ԭ�5���x��uհ�=�(��Y�9�#�*���4�nM��9L�.�$S<�v�^�.�C����؇�x�t��A<n��-��V���g��}�u�Cߝ�z؛����^6�=hGěv8���E\bI�8����X�i�14_�
2���N�����w� cyq��Ĭ�#�O0�^��~p���E1G��=4�8.��k���ÉW�F��"�G���BÕ]�����X� ?�Bd��@�%��<�%�c��-Լ�Kԧea��9�q������;��S�i���:8���H�Ix�6AĚ{��] ���a�=�jMH�0$]�dY�#Dmf��8h�_=vG����p�u9Ǻ�1����S�@��h��=&y�$jN��l$��kua����kE��u> ���.hO�}k���:F��7��F;吝�)����?p�F������NI�й�K)/g�ͼ.��w� ��o M�.�!I�.%���ԶD�&�v~��0��p�B)  �sK�24�W����������z�{�#���TyW���{m �cC��1�	���xm2o-�fB6���A������C{f+��nk�5�5�sKk�`�RT�J	:|#��;��obix��vC��*q{Cn�a���s��:�&@�dk}���|pE�%r�!��Ӥb�������R��a���$6jR�!�{\����F�2�����Y�l�+���ˡ(�M1�atr�7j|�,�'I��0O�@ݪy׊7�w���_BcO$�P�;��ƫg�a����BU�z���F_�r����ۇ�V'�m�Vw��7Xx�\w�c��j��7����/�2�?0Z�w�#�)mf�N%������9�j�+6��,�A#B�d��0�2�����W�Cj��*ECw{�uŔ��8w�R�sB�(�\`���ړ�]գc�X�B`����_P\�K�uM`ܡM�lfҿ��z����$�l~@G*�+Jsѝ�e��	P�e!� $jrI��eQ�&G�x�G\Y�:���YZ�W_�o���#�C	.�P��ò3�Ub�Y>��Լel]��}է�ޞ��m}MgA�V�*o�O�k�}�r�����'f$$���٦���:�~�с��S?9̘gH�z��O�Β@p�@NOy�O:����!n�܄9��-�ζX�ob��R�^et�̳�T>��m.�9+��|ҦWҾ���!�[h>|�##�oݧ�~���z+�sR@O2ɵ��9T'��D1IIػ��|F�=nL�k%`��y��Z*/�σ4��ȏ���f������w����[�l�d��D��8_��Ɂ���MRW�j�<P�A����[0�v�s,g�2M+���G����K�1��sf鍧F1�3ŉN͓ ���P,1_����84#�;gz�@$����8`?
�����/ �q����`܈�|����Z�ݹ(��R��K�����D��#���@J8�����%+E?�I���+�LKlG�IQ�/HD�6�P��g9U��Ժ��]���2L[y&�G*���_�ֿCG���R-����)�� H�x��7��^�=��̒�[�b	�V ]Vy��r�9�+������8�<���/��A�PȘ�j��]�I$͈;33סOU���Z����?t���x��-�� ��cx�}�-k��}����A��o�����ᔁ	���t�kUk
�%��3�v�(3{̂��A�核���i�"3F ��ř֬.X3����۝�ف]�~�_`���&>�``-R���Ol���`w��m��{�{bG�������.�Ӥ��Y��:6HW7���2���]�5H������B�Y��fG��+�WK�x���OQ9UٞT:Zz.���tvbV��:����o �:��H��{���F(����z�[7��>�r��R�Q�i�[�=���k���]�mcN״0�#���b�c�+�=�y����*��������ШF��'�b́&FC��]\�<�Hi��)�R=H��TK�q��Y�磶�m�;�᷍���C̔��R58��g����S�ʮ�q�=`�����˶}&�P[�4 "
~Ӡ2X�%z�G�����)���_+���k��y0̎@��8k�U��蹵n*��-��*�(<|�H�0C�p�Ip�5�J��� d�@��ґ��j�C�?���[e:��Sz�e�S̐��X��nO)Q��YI�c�+T���HI�p�|���;����9'v�Os��kΝ�G*���,���z�qG�T,�#�P��3���K.���|H���O�@��� F�؅Q<%����d�t�����#<�D&_�� `D4�աF
x#�ګ_�֠��]�����G���!���<sWM=�2�����9����m�B�J��Z�nf5����r��
��gͶT�@��:�����H���!J����P��<��-���{��o3��uk�f8�.R_5	(��WY�w;n�_O�G>�'9�Q崵n�N�T(t�H�2�6ٿz�9���I�ˍP���.UZ�D;C�Y;̷;ߍ5�w�Ƞ�NU���h�2�w�S���%�Wʟ.`�Hۚ�GCr�Xu��*�CY,7BO�vԄepaQ�֤���<KgSDe���#BY�̢У��ƪ!�[�|�O6�JԌ����F'm÷��U�3�M�@��D�\��/�{%��>��[u��삑�xPBё�ٱd�����.�e���I���X>�Ź��F:󺚑U���Yt;��d�Sow�$��\F^�0�9�"2�Kr�ܭJ�-/�]�V��j��� ��;�v��T,��GÆm8�� W�j~�&���3.����I�v1s� �k���_&�h��pA��O�B?G��ő�[b�E]�!��λ���$�
�9�1C$�D�D񄩴����q;��#��&����m#QA���5'�\�xz ˍ�+t˧�$J��������b������q���
>P)	"H���]�����Ą����9�s���c�^���^j�����(�� ��&�'�Ⱥ�D�;ڽ�٢�Ҩ�z'�}����`��[����1ޢ�K����B5O��@�X�S�Wu	�Q@�T�Ҕ�.�s��;�(6��u�+����;b�+�Y��ł�g��9�������+�;�J/P���C��ݧ�S��)٘SZK���?b�Z���j=1eݭ:C.����]F�/������b-VJ%�Z�Q0�R5�!�M�+�����������X*��Xm���}�L��aS�T����,�[��4`V���bP͖�ҏ���_�=Yx�M-��װ�d�9��R�;5���I��ױ��i�2	5*C���w��>��J�8�B�ۻm��[�,���2�v��Y0�<��Y������VO��,G�7V��|��js�/�y�&�h�B?G�֙9��qƿ�y��;�!fω�܍�$�uђ���d��f!B�v�1	�cŇ�'�������2�
��Z�i�"��m���O���-��i!�My[��_��Jݮ ֱؘ�������XO��s�WTv�Ʋ�h�lHJ|˕[]���0|Cc	�|�*��%�Y�~�����A�z��"�]bO�_�;-�����A �d�*1��,͑q'��I^�P'�V���V�·G������OΥyQ��2��w�4L��-NU�e��08����ڤ�3ܬ�b�9Ʀ!9��h�ǖz1H�{��_�T:f�C�P����HN��EarI����T0���n1�EUFV~iP�w����GO(��#z�>��]�U���t��N�;�y��B� �LG0L��3]ǅ��%<�c����<Qdƽ�=BL���Lr�%M�j72+xs���"�����\�^����:�ANy�E�^����ȕoM�`ɏ^��!RR)�w���V"�"3 ��YǦ���C�p쫀q<�ٖ�Q�<ln�Rϐ!��ք�(��q�y-1e�wTރ�'T!I���T��h�.e�|=��T�Vd|	�Pe�Q�98��k��ѫ�����K4�٧2�dg�["�O#rm�t�+-V|�kXp�˼��_8�ᩅٿ�%UG��D/�:;�d�(������W���_⼇S�t��u�����1���R�����& 3y/�9�
�ם����~=Wp�08���~�K#��x�����ta���+��?�+�J�;�� &��[�;�!-F��6${Q�b�?`�㪀�Y���31�Ƒ�I1�����A��&1�D��L�n�(���	2'�R��L&a�(R[YĞ%�8Z��RH�
�ѼS����L�2S�P���i�\=��$=�c"6蒫
Ub5^� ��s=*Ħ5�h�?�G\����~:gR���"p��-��E����C]��<l��
R,�
?������sf�d��\�h�z����@��<��K�m�*(��-/?n�:���･�כ@��f��uzzc|3��g���/���&cN�Dr%w�F8#]`���;q���١e��2:��iޯ���\O��9-e?�����L�;Nq�Z����ϕ���HITtto��?�z\�>���E;��P�(k�&\�a9O�!�d3vH=^w�B'�9�.�BN	Qr��T�o�y�{Ѩ$�[+�EX��I����Qi��]��Zg,+��E�t1G�2#;���s�wR�U�J�d�5I0�b6Z�Ҭ�5�ŭ��P	���Wa���1��e:�b&�(
��r9�ǛO2�E���jn�F)R�WI��
��U�<��_&����a���Hy���°�26ϖ�����������z��}��2��Br �U�k~ڂxk'���aG��f��{ڝL�)P����DV�'jX�b_<L^��^�B�fp6�t�_D����5xKP������$dTșc�.\J���.h<D`iS3���^;�D�:]�����.� i'��l���ɯU`����-
��
-���}���~�� �
7Dё�/vX|pƼ_���zI�J�`Gd���(�_KIj����D��{3�jP��Z>�[�	a�Whc3'� 8}FS�Q{��\�?ز���]��.T[7�C��W���9�(�����{.���&�[�ִ�vnˌ�`3%��Z�}tʟ�я�b,���n��X�^��`�As_�~�L�g�?����`�X4��	V�)��ፚ΄�m�抵�����>=ໜIv
V�������:A����9��b\����KHO �;�j�S�	���D�����w��2���2�<�>P��j����7�H:7����h�=����w�u����[l4}�^�w���o=;�H!q!fI<����1�(2*��PA9��/ob��t�;��M�7Zx�z�Kށ]�82�%2���&�Pe��(��u��7�a��6��j�n�tǆ�s5���~�dѫ�8ѳ�W�CD�䓧X�D}��I�f�\Z�����x�w�a�/�цOXS��Ҏ�Z*�k���a,��_[�@ٖ�^�?��!�93	�~e�t��ذ����:�K��Z-y�g�ȹ�ǗE��5�(�HU  �Ĩ��k��y�-�a1-�N��`u+VA�gp�-aș�� �#��l_��a�T5�`u�TgE�0x/�c��YX���c��0��ۡ�$�~6�X�3�i��%l@�?>�=
���~�lC��;�{^�f6x\����nkBD�BA��vU�C�H�4�Ϳ::~h��p�-����0�����uM�H�����3gR���$�Nc>a'L�
Z��1�e=���2a1"��W[e	fb�2����Ѣo:����a�4uz�\4�D����0(��,D]KC�1������$�AY�T�9�Ȥ�,W���v�,�V%E+������������M�����J`d��M�7JP��>W
����J�r�",�0�u�lbv�^�ܒ�0�[�P懲N�79�-�D%S? ��YM{iG�}�_���l!�`��:	pH-t@�|���֟�}�l4I�U�� {�����c�!�I�����u{wS�V�`(�Uu3�z�,�Ii����օ�^���I���6�\���)_,�:���Lʹ	�k�u/M�J|�pEg����OC�5�j��](��`���#L�;gɉ"����Dcϛ5y������י/TL�ʂ0x\G)�)t��y��oEY��	-�K� ��sj��]���ê�J���Aj3(ϛcn��ͪ��ɜ�T@�v�נ�$;����à�jBzPn�,�q����
�Y����
+xw�`k�`B�γ�KH*L�p��,W���� �>�3�h�	o;h�z���3�����vOM}�%?�m����G�`��33�0�*�f��.��6o����1��X��(���{gդH�_NB%T�����z?�a=&fr�^l�C,�y��t�O�.���<g ���z�8�G�iZ���(����=E/��(��p�Z�P�W�[p���4JS�tcB�Y�>�2��-�KX�
_}�=:ca�jwfI%yR��Ǿi�MI�^�j�4L�h�!�x^K����� ����E�8�����<�q+�ԟ��+W'�u����c�A9I�I�pX�o ��l8�o"���UBL��IG��*�(��(��Dj҆�9HQz�堅�A�M��C�!��8��L{���1�O�=�R9S��]��$�)^�ϗ�5�2=}��SO���H:�4�3�m���t"!8"ʅU��F)��H�����MS�V��>!w崲�~��O}H���b�	u�VsGP^:��a��~*�:��ub�*��,� 0"%� ��:Z��%��V7f{���2��ө��?/�>�P��m�&,H������� ���U�4b��
X �uŗ��,�/����؅o  ��e������	7l�=�\��e9�4L���r[��?�Ɨ �^Gc}�22�M��H;~��������{��I(K ������W�x��Q�u���֊˹c�l/��^���e�#��?ۤ+gƄ�BS�`J��	m||��o'��ː�X���LJdT���F�5O�߫�@� ���9�-�G��\���1?!�
���|f���Ā����\&�߈�s�Q8	(�V�y�zN3M��`�6������W�fK��9�7n=���s���T�U:��htY��M�JË��d��z�䄨����`C0	$L�.H��'�C�QZP���*~�6[I5��<��ۖ,G	n�Gx]w#�`�2��_X_��[���$`�U;i�^eb��z��"f9���}���M�iV.J������ڊʬ$��c���bU�	�7�F��h����]ʻx�c��F�����I��yNvky�a�F���̲Y�\h����?Io��l^��!�d�g��5K!�+@M�����P�y7��=ʂ>+�ͧ��
��:�B�ٰДX7;(Ks4&bv���ȅ��K���?d>��t�q���U��7ž�K���PQm��z�Ӏ�]VQ���F���5p;��8�����&X��;�Ոښ�:��sP{��N7���>V�3V���ZK���s2"_���4��T.v�`�J<f��R�*yWK����6r�������(��Pʥ<4�̪����7��Kv�Թ:9������d�SƩ�;�-�����/�.0Տ0O���o�����eT�9�t�zR�d�hl�oz$��丐�_x���^�!0���Z�{��s�9 �>5�ĩu ��y���1��