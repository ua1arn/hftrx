��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-Vț�UM0�JK �73�h�J��ŝ��ܽzAV���.�z�POifK₿7�\���"q�������.p�<H'�=����B���=��t�����!�����\>a!�Vt��@#uG9��P�r�i�ʒ���u�^��/��N���H�ؼ�Ǽ�+���EC��!�ш@<��=3Xz�'��L�E��e��=&�D�=Y�*�H��G㚛6`��r��`��D[�Y> !�o��r[$UXx��t�l퀝=5
X�&�ھ(�;������'|��������� ��Cn+|sy�ac���i&�䱜H� h�G9:�}�F��iدP�S5�\�,�@oFֵ�EX�):�S���P���[�򫞠hh)v[҉W�h h�.j$�tY��4�.�H��z��М1��=V��>?+�~-����C��7)?��<��� cS6�34ʱ%�N7��,�}�OG\5p����E*#_k�Y�0}�GQMN��B.Nb�;�9�͒ۊ�=�W{��3+n�
��VxI�M4�G�Vn�4܃[6�s���)_]8�����x)����lב�@�B�|~���� ���V�!�^ c�A+=W˂���1��٫	n����%A�'�r$�L��z�˂���R`wc<�dB)�4*���22;�)� ��3d2�(db^Ƽ��Qв�7 O���W��A�PF~�w�'���T�y؀#μ&�*P��Dhi���k��p��*��om���&N�Y%L�_ݤE������*��b�4U�I�쯈{<�̀���4"�	(��i�h��t�Tz� Ԋ�L���;`8_´�����X$ڤ�p���}㿯�<ڀP`��E��L�U�D+m{����3���|Zx�k��m
ĳ�g�0���,py^qwt�M���F�´���R���d���4a��bF�6>4���ޛH���)��*W��{1#y��v���'%�����2�=D�X�����H��:J�[�]�녾k5W��YjX47,��Q������#��A�7�����X���7*9=G� H/jH�\Q��q�BtC������VW,��)8@��9�� )Q�C�e�Ҏi)��-8rC��f�hN���f�iY{�|�f�Pc1.ӷ��������yJ�̡]~Ф�L
�1��èH�ۥ+m�؍.e�{B�U��pu�$��1ۺ������8�9LJ�~Z�!�b^�g�ɢ�_@��%_ч�!�(�4^�a�>��Qb�y}��L���A�?~�܅,@�ε�.���z/-��,�~���|/s^���.3�?N� � /A����Hr&>ڨT�n��ҿ�k&����ۧ����cU�	\�FD�뢉(��eI�/K� �t�7}k:�X1ytc;�l�-�
���b�4%dWr��C�q螹�A;w[�J��q�]����J6�yƑd���ԕ�����P_��9�����nDw2��B�L�$�K��	���LбB��}׏	I�=ؿ���e�+�b>����k��?
�~�B��'�t�JC�z�Œ SH�Na�+ׂ��J�	�q^�S?K,W��*^8ݗnq	}x��r"n쥳�н����*�sd��3�0i�Qw�����D>)�=�(���Q�&�4���p3��?{y�x檂���mw��Dhs��:�:�!����:&ByS�#���.L���F�ri۫v�zBC��rq����������B;C�(������$�ͯ�q���hn�R��b}�zr��cU�ށ�q�g���wI��"��.����l|���N[�Nfz��9�:"�v<�ra�'��_e
="#0�R+�<���n��Q��z�#�-F$�e��Ko�΋�*%F<�Y���g�0.L68Qc_Z��v��S�˟����a+zB�
����j�P��fI1�7`�Z�9�9��"vWf��Y`��i#;Ʈb��Kh> �={["�y+���q�?d��j�0(��S`��ܫ�Z9o$=0��]O����F�>����� �I�O`v]���]� �O�
��!�g���B�;N��~�ڑ�{�c�RM�g�I%0.X���N����RR�A+���C��:���9aB�y�ƌ�WDO�D>�.���s4S��u�3�m<$�H�WW�~&��=I��|�f�� ��+s�KI<P����K����yTa�T5n�J�ty��&1��"��$���:NU��<c�.	g,66�5����d�HP����o�i���^��8�e�݌�r'���<U~�wf��d�Ìh*l�xpu�,��Rw0��։AWbȢ�s�4�Dxt�6��, ����}�tj*��#bc9%Cb�Z>�f�G����xf��Ň�?���qM҉*��	��=X[ޮ��PO��e.���}��U$ܘ������߫q��I>�*�xi�;a	�ʥ�U�R1АO"vT>{BJ@n(�jG%ޣApD$�h��^�lS7	7�ms��oV��4"�뮷��x�:��0��ƌY"���G������`%j��	���{{Q��`G	TdZ��+����L��o�#�P�ȳ��є�b��[MbD�@X�a�I���u��&���wJ�b��M���-(6S����R�'����U2��������Id����`��B�V<�����H�����i�v�^�d&�����[��\=��D 
$�sAG�t�U)IuT��-B�SQ\�����W���~h��I�������>g����l��=v[�ϐC�3]k8�7�Cd��w��%�����&��8�`in�M��j����S�(�B�B���0J&��?n��|x��"bA��@�{�#s�<,�ŝ�flwU�h-?������Xxb��ᮦI�o�>��8��7l�����[I��a�d�V��rNݳsE//ұ������ϢH98^i�#��4��ֺ�&iU�*�(�B��u�C�"�O�%v��%ή*_+�y?�po�]j5/Њ�������k�.<v�X��*�t��<�G�"�7pɫ��t�/�2�r�\'�x3��yG-�IV\�#�?��_���4 :�&h���&Ux�wped�&V�+��T�2]4Le!�,ta�;��ND�9{���[��������ΕNkX�ģǰRmd���!t��[둛AAS,�Gïa<��M Qk����|ɩ�2jy��mX�*4k�0��o�n/Ip*v؟��|���,anyMKp�C��J�ۉ��!�=M#aض��;���ٽ9S�W�*m�4{��5{\ks��e��do ��F�l8��W����Wv|	�ơ��R���?+��(Q����S)��_{<A���X.r���)��l�O��SsB~k,.�A�|==�����lZ�4)"'�Iڶ;x����$�7��f�To�|�0�A�����5�{����]�}�:�.,�#��P?+	-BbޒL����.���{Z4��s	G��\��|�q�z=��l�V�1�?U�p��Y���#k!^4��Yl��`J�6��=���i���g����}cUkگ9�����o����\u���[_�k6c��Ѝ��p 2����'�Ş)�d�D��K-��`�<(wŤ�*Q���:�>���hrkv�>"Ps�?��;�L�8���t��j�@Q�	Q�EF�V�X�f��>ߨ�8N��]�%�?6M�J9;i��!��x�2U`z���f�P����JwG�F4@�c2��ƚo'����P4���2Q�`��?�CM[����6��i&�qd��E����Pϐ�
p�W?0mI�n��+źWg(&7(?���B�	U��g�HY��'~,>��.�x>�����<`
� ��J��
G4�����cvh��#�y���C���h ���+�[������ ��?!Q�o��+Bϰ��8>?��L6m��_���@s���CIX�..~ ny�Y1}��2�+ T|�Z�>��ɑ�z��w��.�zu�fLY���<˸�(�H}����owW�Z_�:a���z�m���*<���fG�$>�M&�>�&		�c�+�l��3��cb��-����`��e��8�u�?:�4Jb���6��Z#��`D�'��D�%X{��J����UD0���K��L���
>i��0�&�|8]�&�4����ӆO�zO�&YS��f�m���8ŠO(�c���za��P+D?(9�ED�Uޯ���7�4X�j��A{�s�n�&��?d[�����^t�������K��j�[���������1��n��N���r2��zC��}�YV�uѠ�H�(z��f��b�7�S�D$!��+�r.�@B�k6��/>��1l��"[��^���`� �D����24�+�l��4.͉�錞���  ��oD�*B+���x,-���