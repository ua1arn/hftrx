��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�'Y�L(�K�O�{��?f���ʈ�.�֏Pc\֣�I��B���t��|U|�/֚��LT�E�9��h���$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA����q�HS�b"L]$7!����Y�f��a�Z��Vׇӭ��!�`�(i3h��8�|�g"#~j[O\ڀB��+ H!�`�(i3!�`�(i3�f��)<t>���PF�!�`�(i3A�"̙��2�����Vc2�����Vc.|�('��r�dZ��߉�󆭋;2�����VcЁ=�t�!�`�(i3CS�Y%��t[Ed�+֚L��2�����Vc2�����VcϔJCS��G�d<��2�����VcpNR���b,�ҧ�ɟ"Y|fN�:@��翛Sf�\�_�Ճ܇���'o�fqII��*�T�٥��T��|g�S� -E�7*����q��jlw��JF#�dnE��k~xhd����Cr��1��i�Vw�oM �%���bv.�]ֶO�4D6=���i��p�b�G!��Z%�6�ǀg��i��vp�\��M��ڀK�_�rۈX饿��!��o���ݯ_gWgj"���\r��3ة�K�~�'o����֜,ӘkR� �KF
������:��ۜ������;�Ӏ��B[/'g�`	�K4̓������9(���'�Pw��[#M��*�v}���<�LK���i�[-z�g��hs��%�-h���C}�{�c\dnE��k~xnE�HC+��3K�<�s�������5��w�:j�.Ѵ�����T�'�"�ݥQ����2O��'HY-(�3�(M���O|x�Ͱ��Y$��7\F���r��RL�a))�kc�߇���G�/9'�$���'�r{V.� !�zg�Z�$充�pje;��M͝75#S9��%V��"����ʉr���u��w)�Sl���-�ed�~篟|��d���Y��^"� �/Jџ�_�v%�����:��/�|^��D"���b!��k�8���҆�|n����wH�L��Rl[���.���M�ѕ�����aWfL1�Q�j+�B]g������Ⲕ�u��w)�S�3k:�(�-X�7�j���,Ud8J��$�ƶ��Ÿ?%�b8�<�#�1-@��%��Ձ�k�8���҆�|n���)kd&Z0�i&��a�&����?ʳ�W�%"4����*�T������|�OA�
܊��?Y2���3m�!=�y����h�}D�8����8Y�&�\�#�W��a�erp����N�u���u��Uy�PD4KU7B�����<�[0YY���\�4�sP	�b\qB8Y�&�\�@N��B@��2�o n;�q�m���mi=��B�-x=�WD���4B'���S�K��i|ٓ������v9{�$W
?%x�+�� fג�� y�dH�]��/�2�-�]?�B�nI�4q�Qt!��c��<%>ì�oJ5�%,�k�W��T�٥��T�Sҥ��|E�EYZ/� c��(�U����	x]�<���e��8�t��s*ո{�x�G�F�����OwꅂF�-!d6߿��b��'�� |X��M��"�D�u���lٽ�G��k�8���҆�|n����{y�ڋ�jV%[&��\�۱��ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l�����������f�ئS��.V&��B֥/~.)��3\�R�F*}�c}��uO�Go@3w��0�c��]W�6������qM��D�J����S��������Ǜ�>�xj���+�J��U<o^.K�}�n��&�X&�V�.Ю �{��,��b9���1��]2�?V�Ľ�߉��ə��Q�^�y�zL͊�q��UG�s���q����E©�ʐx�?�'n�^0o�!���!��6�e�:r�"(?�M�_뎱�:L��ҭ�Y�����[�����cJi��2�S�ڬ��M����@qzL͊�q��~���r'�+0�l�R<�q��f�}��h�'f R!�`�(i3c��Et��q���U�ЂDa��(o��0��7�����5	���]���>����C�n��J�
��!�`�(i3c��Et�Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9������>7�,g�YӅ:�v�ј�"��Z鎬�����
��al>���,�۽��E����F��j��\w��0]����jq��Мl�v�ј�"��Z鎬�����	�7 �#�ԬQ���g�z�&����j��\w��0]�o�t���˩��*���]2�y�Z鎬�����	�7 �#�iK�D�b=���>.��j��\w��0]7��u�����a#�fv�ј�"��Z鎬�������(���pl!�6���;b��g��U-�e�,���6+�H�%��ZtV/u9������-��%Mό���.�س���*G��/�p,N�By3��<�]�!��	Ǹ�y85�����3�|#9������q�D���/�p,�]2�y�Z鎬�������(���/��A����Q[R�7�}��C˥�2�6�d�f�����
L'���Xwp�����ʍ�ڑ����E��@IE�U��>��l%i�-�Q�rV�Fg�YӅ:Ԭ����
L'���Xwp����c���i�L�����E��@IE�U����S8�/ #O�)U��֜��3,0=]^	�&|#9����m��
�����\��Fw�]2�y�Z鎬�������(����F�dH�/�R�Ĳ4�������`y�����i�����W��(��"B��$I��w��,c�A�L'Qī�*pY����q�����S�ڬ��MN�ދO�����`y�����i����<)a��/8f�"B��$I��w��,c�A�L'Qī�*pY����q�����S�ڬ��MN�ދO�����`y���C#/<���qg9ۍnJb�
'��(�<��@d�Yt%�)Û4�=w�l��ǐ3����=YN6M�Jv��4�vD�a�ξ���I�2�W� ��iE��G�����(�
t�ژq���U�K͔�����Y�b�Δ;���}�I��w��,>����C��T1�8K��FR��a�z ��(�
t��Y�{'%sAX���	q�KS���K����)��T�\ ��Tǯ�!���\�<�dQ	���qk�ZV"���:��#tCE8�^��㊏')����=.�����b^�'2���hk��&���#�{�0;�}����\�w�Y��k��ı����V���}���s+���JrC��
�־���1�m��P��I��'����cԱn��aМ��IÙ=�H�R����/�R�|_v�:��j��ji���+�z�m_ �e�12Rq�L$�t���1�D\�;b02�O���V���ӕs ��Ӄ�m���VK�4�*�Z�.S����%�z ��y�Κ�9�"�5z���Q��4hz�<Ρ�Jn,���`�rs�i�jf� l��E�4.@�7��y%%��`y����@����gG}O��05GV��#��6�d�٣���N N�S��t�����e6`)K���U�g�q���U�NÍ:��$��fF�:�����,8g5�e`��9����� +��Q]� _ό���.���s6��ݓ��E��*ZV)�J3'T��߷�d�٣��c�A�L'ϸ��%\A�����?,0=]^	�&|#9���b!��u�;s�e�$X�I�K�9f�7s�9���o>��l%i�-ݓ��E�e���F�&΁�a�n���d�٣��c�A�L'Qī�*pY��am��	t?�*|�c��T�\ ��i3�|)sՀ��R�A0^L�ܲ�k?��i%Q,$'���Xw��9�"�5�-ďH�V��#��6�E����FZ鎬�������(����F�dH�/�R�Ĳ4�������`y����@����gGf���3{�&N"3A�NO��Q]� _ό���.�}�
�?��`�mp8V��%�TgR'�n`5�fK��0z�cUL|�]���?.�9$[{^7��y%%��`y����@����gGLǀW3 ^YO�*�q ���Q]� _ό���.Ӹ@����gG��a��� ���(ғ�vq�\[$Q��
�̞��>����� +'������݃�Q[R�75�e`��9c�^[v�5�����N}�d�٣��c�A�L'ϸ��%\A�����?,0=]^	�&|#9���b!��uፘ��|�~�ֈc�S��b�7s�9���o��S8��<�J�QM����2�E~9���i�d�g��U-�e,%�0g���z���Q����by��F�E����FZ鎬����^�d�1�a̳
�CӞDy������!�`�(i3�d�٣��c�A�L'Qī�*pY��am��	t?�*|�c��T�\ ��i3�|)sՀȄ񕲿d7��xg�jзq8�Ј'���Xw�j�7����w�K��ݑ�][H5���8�R�wX���wP-�H1� U�9�q�b��|25�e`��9֯���,s� ��W�d�٣���N N�S�qg2�K?\�T��Z|�$��R�lD�]�!��8�$LQ���qg2�K?\{���Sֈ��]�!��8�$LQ����&Y�j5�!�0�lCR�.S����%�#�ڊ<?@���,D� �6�0Wv���f=�N׏�E�@#�8�
,FIݪ��	XF�t}��oC�H��M񈪔�J8��P`S��|�����Q]� _ό���.�}�
�?���v[2�!�`�(i3�d�٣���N N�S�qg2�K?\�3y��5����'���Xw�j�7��a(􆿳���2����.0��jOT�I\��Y��{�%��^�'���Xw���,D�x ��s+1p�أ�5�n`5�fK�\w��0]b!��uፅUʮ�V(Y�)�ߡ!��]�!����w�Հ��}�a��>�A�IS���2+�R�F�q���U��@����gG�O����o�!�`�(i3�b9����U_�+X�Ă�L�i�I'�QFI�Ne;�z���Q��ì�u"4� ���3�Һ�cY�~�"���ʷ������<G��MyA��u��Y'GMSc�����E����FZ鎬������_�,�;�7���c����}�����Q]� _ό���.�}�
�?��Pۢ����!�`�(i3�d�٣��.���ᣓ͠�cEp	���>P�2-i_��VzFI)�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��_~�TP��b��@�(IM58��,�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U��z�C�f�k��+ƣ�+�ه�ݮ{֯���,A���A�({/$�ߺ��]7�O�e�^���N4��|	�WIA~�R�$+��T�!�˭�<��a�X�c�S��bƨ�_�#��H�߳MkS�QQ5�Ӆ� T���7��f:���t�UW���.S�QQ5��ܲ�k?7��f:���m�
���n�%졿�p�<���d1x�&��Eėe؅��Θie޸XhZ��Q>ml��ݡ��1���I����~u7�UyR�j����r��Py�т6�-�����;qY*�Ld���Q>ml���ʍ���I����~u6�!)z�4�������W��(�׾ŞWsuz'���Xw�j�7������on�b�Bϱ���\�yGL�.~����asߗe�`ޘr��;���	p+J�a$�Y ��!���c�A�L',� *�]���NǨQ�b�ߧ�_ρO#��]��3�u�0��Jn��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���\���3�j���;#� 9�Wv�A���Ibe���W!��T���l�T����ge���I5���!��[���\����#�G6d
�Ld@��c9��EOX$��)܅�����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�O�5�T�'G�+R���o��_�Rv�䩲$���dS@Ɵ�o��èVxjzӝ���I(͂��-����'�)�������9�x�\M����@|����^a�nu4Bޗ��jw�	��x��7��74/�����w�`L��t���Q�5ߧE4��Fr��jL��[��M��qx �i��TpO?E���Y�`��:!
��P�Yh��2gu�Kk���
���/[�ڌ� *�s�ݚ�Н�!�`�(i3湫�5��Ԧ�K��9����ᰎ�+1��<y�3�g���f�,�k]A�|�'���!�`�(i3!�`�(i3�A!�,�'Y�Ҽ~�ƣSiI9�o«IX0F�M��u6%�T�8�w��U��k�nTK��scX{�X!,�0�U,�3��Y$�VZ�ڋ���Y���GiL�~��H�������+1�;�.��1���,:&Ȍ�g�F��6b��<mc�lv0�9l�'����u��r��!�`�(i3��w�`L��^��&vb��}Dq�f���Ě���ž_�F��r�-&�&U�)j�S���ܚ��@��f�\%o���LET;�jmT�#φ��<�6��`䘸�|��JB��]���>���F*a��o��х;'֞�ax�=����h�PI�	mQ��5ߧE4��!�`�(i3/�"����V(pyL0DMlE'�! CH$�I��*�M/*�3��7ݽ��!�`�(i3}�	76�&�|��3��׹��ܜr�a1r8���I����ht��ܜ�[�^���H> �D�9�{*�,6����Z9��J���笺$gQy�f���@Z���OB�n!�`�(i3��7I������\��ʳ�(�^���H> �{`�i�)��|ʡi��!�`�(i3{�d"���e7�[p��2�ϟP���x���^�Q:��T(���27:�������&2��OY��+���C;P!�`�(i3{�d"�����1 `V�(ќ3s����Y�
��<��U�ӿt��)"&�v�"ǉ�t������z���!*��*8�N�Cٺ��#o�]�ʄǡC�o��vr5�Dѯ�e3J������f=�N74/�����[��o}��MX�w����D����K�f��9Ƞ��Ծ �����]3��>�O�i@5*��^H\�r�� WF��=���Q[��>�8���q�p��7YB���@V�y$wV�I�j�ځD��d�N�d@�>/�LA7g�
H��,А�r�fDT[Ϧ�31�"]�Y@���.�%�{yܾc����o�&7;h����*L¦+DS�%-4o��Iuu��w1j�Q��i�8�F��(�[�o��_�Rv�䩲$���dS@Ɵ�o��èVxjzӝ���I(͂��-����;�~��-�f����Ga��'DV���b�z'hۉ)��d�7�qĮ̢k���F�KD�Vr[/}>5��0�B� �b���H��������]��	-:ba��O�^V��q��� h�ҩ�7��u������v����?��۳lU`7�X��=�$f��_Ub��7��G_���;�P�t�5�׹�4��)'���-�5k\u�'A�뀉x��[�U�\`���!���y�a�����o�u�/p�4YMD#��aՑN6h>���Q'i�q��p�u9� ȫ^��.�')V�E�L��N�?��~g�����%铿7@c���K�(e��V�Nyw��aߪ��;̠�z��!�pF�?�~���D$�ώe�LcQb/[��l�,��Sǿ��U�|5 @H�/��z0��j
��r`I��4��IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��yЕd�tuљ�FdG@dN�<@Iv��nt=:��:5A��p���N4�@�S?�Pm�/��kOT*qA����6\�4�@�� �-j�1tSjv�F�6�_���3i���Y�
��<��N�g�c�`!�`�(i3�W�3�-����⣮`4hz�<ΡW���b�0���������5)��Z^�h��N�M�ob�H���T�ì���������;b�-�2��"橝[��ԬQ����5��t�	���QC�꠼*d�m�d��-��!�"ǉ�t�0/0`9N1�N�g�c�`!�`�(i3�W�3�-����⣮`��+�T[n�����$�~�+yp�l���d�L������.��U)�~[��Q,��:5A��p��jVѭ@�����$�~�+yp�l�#QSU:�����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�qb�V�_2��Z��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���b�A�_HyN#"�c]=Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hL�6��P_qk�Q��R�φ��<�6�@a� ��fFMqlg{y����i�q,?5qřy�m��^x=m�� xjzӝ���I(͂��-����>�Q�c6��=�ڹ&��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��Ư�ճ�%6�E~�{_8�Y��=�}�Vݨ��}Dq�f�?��LST�ed9��a��o���H�RtV�^�Ư�ճ�%6�E~*�k���-�@�,{n8_�=@'ѥ��Yn3%yaJ�����ӹ�Z<��A!��-�����d�tuѽ3y��vjLo��-FZ� d�!y�b�G2�Ra])n#2�A����(�w}� z�P��1tSjv���������O=�W���˙�6Ï�9��D�y{~,�H�͛�HN��R��F F�E̠���F��O�\E�W��4b��os�鮊���4cn[ۮ]��E���AS��0+K���t�T��?E-h��`f���sd�G}%����3f��$�uGci���{2�'ž1�|�'����u��r��$����}W �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^����,����0�|섃Va�ir[��l�,t���H[W?!\���k���%�8_�mS8<�n�ݚ�Н��&��>�'�^�����;b�-�2��;�P�t�5�H�������+1�;�.��1��!*��*8��!�qgy�`��vN���+A���o��<�����	G0��t�UW���.Ir��͕� h�ҩΞ �@[�鋽C�H�CW���|e"���F��O�}�	76�&�� Ӗ�t$�)�vxj�y��j}���*��>Dj9�J?�����A"�S	��1�3�����+�}�`��:Ŷĺ��}x4�Pe�I\��Y�tM��楱�o��_�Rv�䩲$��8��I�:Fa�7���z��O��߿�wW��@?��WA(�c���_G��Hb� h�ҩ�`&c�'N�j��O|���/��kOT*qA����6\�4�@�� �-j�1tSjv�œ&|�9�n��~��4�)P<�ܓ�Y�H�������+1�;�.��1��r5�I��d�n�{ .p�a�	�Z�������>w��-����Dw\���I\��Y���*�f;��}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ-�+���5��o��~�Q��g�0��=�e
B�a�\��{3�5���l����#fQ��=�{-��ō܈��VtM��楱�o��_�Rv�䩲$��8��I�:Fa�7���z��O������������a��r$ɓǃl[�Ƶ�1tSjv�œ&|�9�n�o&uL�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b�Ѐ�(���0�l{�]&"(�q9+t�}�|#HK�� ��5%q���f�e�!\���x�sl��gVdxQ,#�%+V��tP"G�wk���zܳX�P��%�©��-/a8V�Ո�����������4Yz����|e"���F��O�}�	76�&�� Ӗ�t$�)�vx�m`���ZXH�7wS��h\K�5~�Uʮ�V(YZ��*x���`�p�*X"���փ��m��r��$�0I&��Ϻ��S����=�Uʮ�V(Y��a��R���t�T��?E-h��`f���sd�G}%����3f���L�yE�:�.�N�������a��r$ɓǃl[�Ƶ�1tSjv�ըa��9�(�w}�W �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�Uʮ�V(Y�t���1�g)P<�ܓ�Y�H�������+1�;�.��1��r5�I��d03�� <Ia�	�Z���q�ZD��,AԢ�a\�2}$#h6��8{4����g��-�����a�}�$�᢯��0����$�a���NM���$f��_Ub��7��G_���;�P�t�5�׹�
r�	O)�A�IS��,�د$�,��B�quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7��vo�V�2�~ڦ'ž1�|�'����u��r��,��B�K� |�>��̢k���F�KD�Vr[/}>5��0�B� �b���H�������+1�;�.��1��!*��*8��!�qgy�`��vN1tSjv��H����Lq�\[s!(���27:�������&2��OY��t�)���!�`�(i35i�a�vb�9�ڟ,AX3�ԝ��R��1tSjv�����l��.���C	���'�PD��	��x��ݚ�Н�ٮOS���p�߈.m��B)X!�>P�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��H���*o'/�Ja�DF��(�[�o��_�Rv�䩲$��8��I�:Fa�7��׏�������u��0C�r$ɓǃl[�Ƶ�1tSjv�9O�m96��\��;�,*qA����6\�4�@�� �-j�1tSjv�-��)'�T��Z|�y�`��vN1tSjv��H����oM2l��Eߝ�b�Bϱ��>1J���wʽqlbך�-����!�`�(i3����@z\��}Dq�f������!�`�(i3�j<��?)X!�>P�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��|`�!f¹o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc|B'o8�R'��o�Qy�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����Ι�e�yrJ�e��8)��0�o��_�Rv�䩲$���dS@Ɵ�o��èVxjzӝ���I(͂��-����3tI�AnM&N"3A�NOE�g�������(ӈ���m�r����t/����>�V��#��6k���������|e"�`�mp8V��%�TgR'E�g�������(ӈ���m�r��������Q��>%L.�A,k������8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�D'm�����Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ�v�4�?zmy�`��vN1tSjv�Z��JP��V��#��6�I����~u�F�{���!�`�(i3�?L1��	���z�Ji���M#�rYӗ��_�Írs��ʟ�r-�T-Ki�\�����Y,�֮����l�鵈R#�K�|TH��A>%�}שĭ{l�,��HN��R��bP�63Z�t�5ߧE4��\E�W��4b����A����q;�4�\����t�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��z��w���0��C�h�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcug7N�RL��{��� φ��<�6�@a� ��fFMqlg��èVxjzӝ���I(͂��-�����9lD��XH�|ը�K�QdN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�D'm�����Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s�l\�=�]y�����ʄ_1tSjv�K��ft���-:��;��ч4H��&��;�T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH�|ը�K�Q5����{�q��Ɨs$f��_Ub��7��G_���;�P�t�5�׹�y���3w�9�ᾓ'�f�
����dCn:�l�U��)���Y;e�iK!���d.��$�Qu�G���z銨���`!'���Xw�j�7����w�K��ݑ�][H5���8�R�wX��d=��¾ȼ\���F�`yx�>�+X�M?��y��M;<QA�"�pM�00_��nF���<�W�.�P�	��
�Q�}�1�:v�!�ӛu.�A�e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�m���>#o�]�ʄ�M��,����q���f�e�x��w����֯���,mk��L���n��<f�`u0�F��a�';��#j�ݚ�Н���c���L�\����<M?��y�!�`�(i3?�8��3����j�4�f^2��ʹ�q�T�c�$�����#oM���a$�//��kOTV�Ո��)��<z�1&k@C�Ɨ0z�cUL��ddՅ<T<��A�g�wɪ��o��:ϱ�՝� s�#���k$ ��YeԿf��&-Q��5�y�����ݚ�Н�>�H��-���vP8Z鎬�������(����.��$��H D��cZ�J��1Җ�u��}Dq�f���Ě�����}Dq�f�ܢץ_�_l�0�lCR�iY�{u��r��Jo���j�"Iե��G��Hb� h�ҩ���YeԿf��&-Q��������M�7��<��am��	t�O8��4a(􆿳���ʮ�����|e"�c ��4�-+��.���!���c�A�L'�ɻ�}?s��{�2V���ś���k��	��x��ݚ�Н��B*�0��IT�q��]7�Zg�x����}Dq�f�"�a�BOPj�+*7u`��]�!��	Ǹ�y85��X��I�ՠHu��0 H��B�%V���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx���$4gozq<����Re��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!$W�j v�'���H}�@v���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h;�ƽ�/����zN�S���t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��y�P#+_]ݱ�m�
���nGW�:!�E�/��kOT*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t�	���QC�꠼*d�m�d��-��!�"ǉ�t�0/0`9N1��-����P#+_]ݱ�m�
���nGW�:!�E�.g"UƄ3[�g�DPp��k��^�1��[��o}��MX�w����D����K�f�1tSjv�K��ft����Y�b���v�Ѭ�����R#�K�|y:�1^0lfHN��R��bP�63Z�t�5ߧE4��Fr��j#k
z��k�m�
���nx�]l�i6�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl����::R�{�>����t2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������h}�"+�{z���K�h�&~pƹR�"J�;����g��徐�ߑ�Km�?0c���<�<��(�;�n _��{�5�Y�w��i9h��W� c�.[K��m��S&ϊH��c�쭄]���Ske޸XhZ[�}Q�9�ַ���5�����,p�ն��95�2����Z�׭ �k�30: ��q�[���1x�"�Ag����<v�Y\`O.C�x��7��c�^[v�5�Z�|��w(K7͍��|��W&":�@��v{�G`,9�H�W��-���֪�K�;˞H���@���4�c[2����ZqJ*A&-�Ri�H����JAA4i1�*_k�B�a��� h�ҩ��H����ڻ�+���i��ċ�!1tSjv�!�`�(i3
/���p\"�!˥���KS����<;�$��У2=E���3	�o�{,\�0+sJ���|e"fĉ>99��A0ok�Ra])n#���r�����Jo���j� ��7P��'����u��r��!�`�(i3����Y̀�3#O�2�B���s�����X�X���`��,n��뾦�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�fF�5.]���E�i�m}6߸��S�Ȍ��9�ڮW;��|Bΐߧ �l�}!�#�bX�h��M���`��&0���Q��Ӏ�FQ
П�мBAϭ!�����D)���w=�ֶJ��:���鄖	~r��kh,�!��-5�M��f���'����Ջ<��0���h*-�#�`���O�φ��<�6�WN줔)8�7�o��;��èV㣅Dy�'0: ��q�;&=7�kJb�z'hۉ)��d�7�q�5�����}Y�u�U���2�B���s���EG����'g`$�Y/!���La�2U�5;����Yk��]�Q�&��H'o�a8��v��ONH!�`�(i3�\!�U�����������[���-����!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H�f�#��(�D�"��ӌ�r!�`�(i3�5ߧE4��!�`�(i31���~����l��Ht5�=�5�G����V/ G��Hb� h�ҩι�+�t2�c�^[v�5�ܾ��mk�9$[{^+#y㪁��i�u״$(�>g�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�Ct�w#��@}�	76�&�φ��<�6�aT��3G?�d���&���TtU��
g1�MVjg[:%w�&/.����#�>�n���X��RLT��T�٥��T��Z��J�~����p�q��l0����Y�)en7�F��(�[�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb� h�ҩ��T1�8K��}!�#�bs��>H�,b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vN�[���}��4N�J�ף������&G�B�'��a��*ZV)�J3'T��߷j��
��e޸XhZ��}Dq�f�m��;���1&��*�("��X2��4�j:��e+�������� h�ҩ��m��
��0: ��q��%��j��e޸XhZb	�fƏ���%>�rGO�D mWN`���*1���F��O�\E�W��4b����A��c�^[v�58u��\B��U<2+#2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�*I��A�*u�>cC=V�g`P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc`��P���P�L29:(�U�E�0�IDKO��	h�{��-�wXB`d����3�#quA0�e�&=u������FmvU����èVʲ��U�4�a޵��	dN�<@Iv��nt=:���2]���`,9�H�W�0��K�[̞��>����� +"�*aPV�6�����Q�8�w�[���:=r��Ɉ�?����2���-/a8����l��Ht5�=�5����������&G!�`�(i3��	~r��k�%�D����MxOܳ����|e"��w�w:�!�`�(i3ʲ��U�4f�
"_��P��]�/F�ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6�E`����Fr��jϤ�LǀN���)��%A���h����u|�
�xr�{���г��r ��T���yo��5�I�B4�٫IX0F�MV�ҁGG%4vkz����`���φ��<�6���w���c�ShT���A(�c���_G��Hb� h�ҩ��W� ��iE��h�{:m��b+}y[�k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1��!*��*8��!�qgy�`��vN�[���}��4N�J�ף������&G�B�'��a����w�蓺���pJ5�!����;b�-�2��z*	��y��R�o�"c�Pd�BR�~;�A*8k��.ͥ�H�RtV�^�<��a�X�r��ڵ�r��@eM�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b�[�؟�-��@뀗2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������y�$��_,�����{S�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc7=�� C7<;< }>�5��Z)l�<#l=��,�W�8"M�5�O�%E#PMQ���0f�Ϡ�����b+}y[����,�ǰ	M,��rER��KaP�X��OV�s���e�58:	�eL�V�l�>@>�~;��|B^VE��P!|�u�ݪG�B�	z�W��7�3Z��ȍ�c�`��H�I����*��	^����-�P����C��CFv$��M�{�|L��ʾ>F��d��-��!g��J�s����0�|섃Va�irH�%��ZtV^�,�/Bh�՘����;�M��f���5��q�P"G�wk���zܳX9�Ϙ��.S�M�#0F!��D�����k$ !�`�(i3V[B�5�mw�R���y>��yС �ݻ)�9�yaT��z��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc0l)�┗u����p����t�T��?E-h��`f���sd�G}%����3fX�?���'�V�2�~ڦ'ž1�|�'����u��r����~Щ�n��뾦��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#���N4�>y�pA��M?��y�!�`�(i3�	�%1A��b+}y[HN��R��bP�63Z�t�5ߧE4��Fr��j�p���"[(�i�x�n��{"[)�`����ǆ�S���Q=-C ��U�