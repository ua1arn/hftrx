��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!����� �@��ތ~4�Q��]�����̆dþj" k�SȒ�rQ4f� 8�$0b�td�y֚+&X�,�3�;X�y��P��Ҥ�,2���(u���4:'�ܸ57+`e�b<g�襧7$��t��ef*�(0�px�%Jc�U�� ���WT;*�E�M
��ҿ�n�-�_�Q���j��i3���j�LK�$���f#��t���$�>�s�����JJa�W~�&I���uW�r5��bӲ�Ys?��k��M�D!�1rP�P��Om�폡E?q ���+G�2�o������L<^W�.k��!߶�E�C[S"i��'J��}�2���{~�DT���;A �0�u7�Pn�I���j>����9�D>���e+K#9gK��N:����ʭ�w����5��}	�s��t#Oi��{�!eyl~�r��͸�Ł�5��E�A����?��W��It����Lz#�[�g`��h�e��� ��T���`�;����_?�+�Kg�;\�W�;����uz��2x����}dO�nP�L(���,D�Ϡ��g����P^+�#��V�\}Jb���,9��A/�s4O���l}�+�ڨ��G
I5:������+?�����|���xk���6c�Bw &ܣq������/�KRB�&=a��t8�{�HH͑�\�R�s?��f#�}�����0���QX�~.D���h�-�h�ԍ��Wi�F�ԝ�Y���TQ%�v���e�H⚕����K������%���dX��=���h�D5GGA��.��j�����3�i��f�4�vu�1b׺-��ڤv�!x/��~�5kQ(����	����i{7 �-���Q���3q�R����[�n�qo6��'Ҍ�^��>������=5��bJ]_u�k�d�:�L����/�Ień�/s�;�J�D��2�<��F�T��5gQ�W���P9��%�Y�5�[I��C�=v�#R-�m�%(;���B�r�G!�iD~��ep��4ϜN�Y��y���>0�#�S�>E�[!V��w{ʹSC�p���u=��E��MF�K�?�Ϫ�s��8�reu�{ȳ��m�>ݩ��kY��5f�UW�y�����^�j����*�Naf�~�v��7���=N�c9"'���X	��t�-���~ޮ8��c`f5�L�U�����S�82L7�]���?��O�ӦB)"2���Q4�2��Kn���Y��)X�ƫl���6��:Z���H�àL�$2� �\�8�\��w%�>�R��+%,�k�/�nP���曞�@�M�lx�|Jf�������]�ׁs���;��s�~m�'ڎ���=[��v�-ܠ3=D�&��h<zլ�K�r� I�ʎ���齱�ˎN6S�_U��s���Ԫ�ѿ��he���J�y�aSF��4��)��G�
��x]����( :Tx'���Ap�����r�Xر�1���]��C�C`����
�م7ZQ�I�x��GJ�+���̕�E(�����70�{CN8]-!ùi.)��#\��|��ap��)f�g��%��7i�Q�p[��,�	���r�w�RK[հԟ/�(L��l��aeO��I�❽;@R�q��Z�>�Q?:���(��
v�4���F�x_!�&N�O@����[�w�7
�
�BJ6@�`f�V�W�e�ּ�#Y�"����h)M�\>?��!cm�Sa��E�k��&
��Ln�V؏�FR�Z��c��"�Sa
���oϫES��v�`&P�WRq�u��1xl��o� T@8�	�E�:LO�[�I\~e�V��I��� h�T<����ه�V��9�A�&/�Ps�f�ά�D��7�4��7��D�Q�?�|N��H��O�3ԗ��b 34s4��BL
*�����$���~[%Y_"I��{�GQ�}���I�k�Z8/w [3�>�M/��fZ�j��;�^S-��_,����"B-o�,���������I��uw�:�v�-�L旋ô��l�[��8�o��ա7��Z'�i�*��Ǜ��̯c�N;�+�R����H�sb��MА!{҆���Z�-K�B��]���9�.�hr�&�F�� ӛ׬k���Q���k'�P��lP���0��Q`9��(����a%�/��������.�Ը%	ϊI)H?�XB���ς�߮/�`�M$<���fC�G���t�7ξ����T������CA����61#�[-�D���?��o�ri���\�R��H�6Ђ{�_�5_��� M��;�3ng��c���ld����x��F`����A�_SWM��cҪ�l#����T����z����S7�ðrWI6j;� �-����MH�]���أI�1�;����;�Q�����9ړڢ
r�Ye���D?��B�^A�O ��.飹�������/�ٛ?�̑�3Z��X1����ߒ������ @E&'��5'>�|n-ݩm6��k�8���!�v��V��(�;y(!�c[x��.ڭu�X02/��:�`�����5& �UT��Jſ؄B��"|�Ě�0m�/�wh���<��``��m�.ܐ$�vm*@���8�[���aO)�=�Q��aD��ON58p���զv��4���,o��v ��^z�U��X�n9�%]`1i�,G&P��@R~rE8�,����Y�m	�f��yoTL�iJ��9��m>~�K�Ϊ��O��S�0B���g�<*dB���J��l����/}<��P@S_�%T9M|xg�T�K܏o�� �Y���}$�������y�J�ɨ)y���_FSK*㬉81C�k*6�����ĳ�T��d����r:��թ���aMc��3�B�Q�Va�*�.��5���������k���]׷��'F��0Л(9��#�u�MS�su�$v�����T�Y�Em[�E�"��W��vfp�-������9E|�0�_�u"ߎ�)����Ʌ� �f|�����B������[hB&8�+�����5qd��<t�ˀUdp���~�hc�����D�f!1���o%�P�Mg#hG���S��>=.�
���[V�8@�O��� K�.��s�ve%���&Kg(�&A�E���V�z��q�� �:�@�?D`<á��xbF�rB���+3>�� �ɥ���c������zb&Α�!-y J#&�n�ڸg��)'mH�K_�wR������5�0�8����;~S\&}����4ev�h-���`s�A�|ɗHֳE��X��
��*P
�A7��jR��`xev-h�������`��%��]�����"~o(.�H�^i0.�k��zP<�&$�όI��@t[�n}n*2�_c �	Ӗ�Z3}~�[7*D�i�l8�h �� �խ��+���l�"��sD\#��9�%�Ng�����7�^Q���͏�a<i==�����۾���[�o�Ϛ��E���MI�l��r�e�A��6氿�~�F��R�L!!��C>s���4���n���9�)��%o���o�n3�[��(��D�t�m+%H���n7�n�G9Lq��I�~X!N������߀� �Y�(u*W�!�1�m��gЫ�����E�R�_�SE_th��#���)����d���n�=ף�y��T,��t�j_��+���2��.�7�P'�%�Rw��c�pK�R�1ü�3��v�����d���H7=n��<�j��p%}~�-�t� ��e�Z~�b�J��?�A��C� �`D��G�W�$-D3�AC�p_ULX�8W���I�H`�\+`6���@������9֩ձE�T������@�Y`���Ҁ�//��[p&V<Y i�M���V��J
�^��	M1&t���'zR�i�`zm�s٭;TsZ_��%��C�"��Z�JO�?��fr��D-�r���C8��0�� �Jd��ɤ�\K�d:��s�^FM�:�:��&����G��LDE;�t錄`GZ!4�QM�^��:U�&��3tF�f/�	��p^��)2ǂ��4�&�F�Z~���"P7�[(�n:1����r\ q�⟊���W.� ��f��W�;Dwk��NMĴd�!�0lG��G`��rN�F��_QJ��5US�kB׏���p�R�Gn���]�e?��Q`UȵD�̤:�����;�o�2�{�4��$߮���q� 2�Zw�W�U�������Zel�ԸE� �u<F��^�s^d�R���5���ʑ�#�L�Cg$(�e�z���o�������xuf�N"�*��_�*�+&Ԯ�1��L�L5�oJ�̷`T7��Ed���7G=ɂ�,lE��P���@�9�{�	u$]Mn�+����5�pܰ��tR�Z��|�Z��!5�:�6���8�������R�vB���ܼ�G�� 0Hq��ױ�󕇼����)����Mˢ��ؐ7Q�9�����Y}�&�
�H�)�Q��Lv�OA~����9�L�Pt<�æb����7:�ͪ%>I���*9�C��@` �RB�'m�>�o]��P�c�O�4,�����g7���sG���=$��ǫF��MR��3C�ߠ��,�q����	�*~�X�v�۾bc^_\�uhC�hG:7+��Z͞���w��C�x�ڴ?8��Z����TJ(��9Pi�\ѦAow��n��V�����ޘ'{Ҁ��l_~_���{�˦劢.*/Գ�8�3���j�l9O��j�@�%�|�&>Q����c)�I�S�$������wR�|���é�uP"Z���km7�f���>J,�RL�u��k�,u~�t�S:�#�]����l=1%��/��'��B]�p0��%�k�z% ^UZ��GaV6���3��ؼm
�C"��	��:5�����I��.&?�a��t��an|��:5ڛ}NH���=P���a>z�B�oX�v�H���B�5^�˴Q��r�n�q��= p!߮�J��Yq�PN>�|��F�wO�ς��l�4�Mb0E��<����U�Ĺ���[u�9��a#��Gg�m�9!?*�G�o��k�؂�q�}�[aW��{��U�5�E�AY�܏ }:� �a�����\e�as�L����ي�@�"|	@`�PL2M8fjRƶ�U�zqFu�?�¨Ӑ�s�"��m�{�w����_@����AU���p�Ώ
^�쥍���l#T�q���L'j k����qQ��e�����Tಹc��矏�P�T16��!u6��l��U��A��}���H�t��$
H1�?�h=����I����~So�Q�^��3>������$m�#e�V1t�*K�_�`uPɵϐ:Oٴ�
iv�+z|�hY�2ԻM'��0�H/�4����3g�^����!*
�/_�+��	�^�����J�W ӿ6���oFB56���I?���_Y�8`h�a�z�}?�ZWꥌ�6��s�t��\:���1�dѣ!�ן��ϰH���Hx��&�'�8�V�I���c#�����3�ٵô�$���&�x��~��n�y�4�Q ��C�э9$s9�	�q&��1��z���)�ʤ�NuQrn�p7����s"�^&aY*��ZY�7��0gD	���p5`򠁸*ʍ ̤�'��E�n�?'/�N���&�C�C[U�C�)����g�x�\�N�ɅH	j�Zg���ł�£��������nYq���V��82�&�qC�3�qE�9&2I� �����\0���@�I�Lm���d#��D��oX���L1J2U��. ��4.�%�z�G�K>i�4���%6ꅤ���3n��8���|U��J�f[��o�%�D����H��a5с,z.�ѷ0D�O%U.J�]�6|�ߊȔ�!�0��N1i�42�lt*�_���*��b(*��ޢ_,��<����(�����ȏ�"���?����63��s���7�y�:�D�u,�l~V+��_�d`��u�,�z�og��1#-B�Rn�G���q���,Ȁ֝�cx9c�!�g0�f�Ė8pL~�͒��K����eC����D�}J�9�]�e+�:��a�!�&�1C��������5&�;�O�l�7�t�HW���c�yy3C��FD�Z:\��(2�c��Q�������4�A�duT"�O� �Ȫi��.�
Jv�W[��F	E���x#N@ |DmN�d�O�לc�����?)��ʃH�ܐ����	g4�Q�km��Hnu�b�C��ތ}G�8Q<:P��A��R?�*�ԨbԉU3Y��ӑ�e��#�4�?@rw�ʎ�|��ѵ]������+ho�"1��EC�ݹe��1����4����2�9VŰ#J�U$��V��%K�B;�kl�Gy��c�G��e}��#rg�6����w��' �&3�{�`b: ��<�F��ߡ��b3�RJ��M�	7�}�4ډf�H�
d\O�<4�D�M�E)i��L�U����-y�xz��������Bb�����%�Kr���b i���$^x�7g�����n���D�T ��C���g�'���n�
��0!���YQD�:�G��*|���o��ղ"�]P�琙��5��]aN1���F�yt��5 ��V�b����pm~O���[�����tH0�=%p��?��S�q�$~[Q�F��C^�N�����%I��h*w�$������{Cǅ!��0y���P$�D��OJ%̡?��G��ZǊ"���F �9�'b�� h�r|�?F_Z�i�{��:�W��pI����A�{@��6AC�#ٰP�>��Z�"zH�z��Gv8%��/���`����3����S �h*פ3D��c
�z���T���v�o� �֩x̈́J����H��	���Q�~�&\����I�4@�`�;S��
�@���9�/��:�p�,�AQ�����,s?��Ռ�<Q__�ʁ�u�
����`m5?�	��+�����6�V�f���
,�LM��^s�0���vՍ��n5oSF�.��u��G�P�"�Cv9�Z��w���EM���d�x:�b�rw���_���`裸�æZf ����P㵻��o����]�F�Q ��E��}+�4�d��H�:�U�Ä2*��~	�g�X��6RG����D�n� �,2�na����'�ȏp�����}"��U���^q���q97���1�j��`o���݇Io3c�g�aW�K���9]�¼�ߧ\��Je�b};8<Ȋd1�De����&#0��P�S�#}6� �3*ƟB�m]Һ-�_�ͩq�o�_ f�²�MX�{;(uB�Kk
�J2��K ��)�8;z��h�(�@8�Ɖ��Ѕ��׵͠g�
7ڷz-W�&�c'����i1u�)W	����7.�#�kT��	-K�)@�f�4ŉb\��_��Y�J�: ne��0�,�8/���>�c��wl��Z�%�����C{\���3g'y48��P��F�q�|��k�A1h���h��)y'�>����{�9#GSbj���{v�P�'��C_��D
%��6�äm�:hϤHDT�LG�u��	���^������Ͼ|�����i�]Np�M��Gj^3B;O2�\U�������Ԧ��v/���)�y���̽Qy3&�vZ���"e�Z����T��T��u�c�7}=j��ff�3	�ϭ�w�>drA��B�]��|۹u.�/i���72�ĩ<�ww*츰Kն{wL�p�ˇo]�,�T*��7׵>�k�	�ԁb�.	�~".о�I�}I܋.�M�%ө����J�#�9�ӕ��UG <�[��o����p�؟`=���l�^��œ�3C��=�\�#��a!��BM�l�W�e�	��" �동��l{�=i��EVIgp�)�Lh�|Ϙ�k>��+��LY�j��m<oN�$c!_�hDz�g�6����п5&��\�]�H�_����cx+�KH?(�}�F��a����P!2[ሒ�lOj��+��Q4`<�����Y�������'��EE"˂�y�B��+�y�����x��
��� �m!!>�Xd�Mۻ�;.��3�3&�����귖Zi�u��6���;ؗs�E�?v��`Ź/"K�([����ϩs����������~[��>���,"%�*�@���$��h�Q�.�8���k��]�2�AR�6 �s����^�:z>���2Y�?Eq�E�_���o��H����SԳ���t����KC����b�6�p��l�����x���4������iAm�\!13*����1dB�m���Qj[S����=03��I�!<��V�j�ϯè4 �#��沴�E)��i���	��[x��A�?U]%.�!Gȋ!F���&0��M�9��vLz��/D �KlJ,2�U�pm�m�gƫ	 �Wz��sI�'٫=#��僶������K}�8Ʊ�+�!4��Q2�������GQoq�Ǧѹ���ej!b��{��D.��������N���Q�?�/i����T+���ǅ����:��x�<1˥�U��BЯ��?X�@�+�����E�E�b|m����<�����1����)�怮�O�9��=�#ߜ�.�="3�8ٵ��KaI ���JB�^�<|�k�i<D�5m�ɝ�y>�Qv�!э��~[��Ó׸K	^j�d��ˊor`�Lū���f���iŲ�Lq�!{aѨ܊y�:�V�|�X �P���Ըͼ�9.���&&$�H$)/(�-���A럸�����@���ء�u���J�MM�9gT�=34�u���)4t���Gtl�٥2���F�en�7�&%��HA�S��H^�vL�`'HС/�����k�1���I����tKE�
�3��{L���%v;���r~-�(�ߤt(*<��x���n)��I_�v]ȡ�=�&����0�nÖ򈁑(8�gL��\�^�}��BJ�	=l�A�ɼ���V��F�8E�yWW2����vV]i�}����5����'�\m�RA/(�1�&��#4�L�a��6$��a�����&�粟CN^�g"���@�P6"K����'���p����P5�h
(5|���D\Q��F���|OP���0��WW�F���d�U���{K��g/�lw��f�ٴ�1�J���� I�8�ńh�W!S��?m��%�;����BsH���/����C	_�h5�<w��O��>��j�u5^<�K?F�12�����%Pe?��V�X��	pC��R�8�5�p�@vr^���C	3�Ή�6% �F�yK��zj��]�Ն̼MNU�Ȥ�q���s����׮���WN/��lL�_qǶ���]��c:�a�j��-f��ΫF�d�d�����l�+�kQ�y���W_X�7�G(��;�V��L\�'���Ǯ��R�{A�o�`d�o-�뙲z�:{h����*T
�S��LLvU%����ǵ���
(x �ۢO]�����e�R< e60��Ng}�}
��5
c����C���gҮ���fu�С0t�RT�敡��E-\8X~���7���S͖,�*2�z�@��=��|�a~X�)&'��7��kۘ�u����� �ch�r��(�҅�dk8I!'������)�
P�,&f�2LI6$�H,���25��:
k���ў�� ���W�*��td�m������l	j�8���v��Y2*����h��Iv�$\[�ƧDo����/!��ƌ*�qb}�y��Sf��n�S ��-+��)�l=7�����5���R�����3�dL��D�o����kG�b�w��#x�$�pԱ.0�jU�a��7p/��U�_=�aMF�/ג�J���~mm3[B��ݐFe+���&����±c�.Y
���!�9��Ǎ�"׋�~��ϣȢѪ����^����sJN��]��˪�q��J���2�M_�,o���!����� &�����q��� 1���e��{��O�s�r�(Q� y�M�ڦ���D[�鈘���?�Ƭvp��
uj5��'��&���<&+���Te�
eV�ݺV��~�#:c>s��A3��>:�b�$w�M�\J%>���_���<�%�;Z�?��Jd���0$ޣ��#K��9.�{k�~��.o��)�jF{���5��$�<\=%���t{����12��k��wh5��"�?��(I}�,[W(D1�L`U��o8v�E����ꔌ���W�і�`���G�FLI;X3@B�����|cO���I�������@}��A"�!�:���������-��yh�����Q#�;YD�Et�zp���s�|l��}C=���Jb0��ĕOSEzvr���ڧq�O���6�
CXi-���[Y���p)c۳A�ڞ��N����Uy���*Ǹ7�Sg�k*���G+���~UD��Ŧ�K.��d*��d�ܨn"VW(F"S29�a1�}
X�x�j�:�*>2n�F��	|r�zQ��
�演���\ۢ��P�Z]_.|�##�ϬU��Za��g��ߥ�t%��":=E�6���Vv���A��7�
���$��/���-�������I��'�k- �O졽�F?P� v��h�C�v�^2'�>� K�J^�����.O}���X���A�O�E�-�)�$$΂�
OIx_@ ��!�{5!����-9o��L4(X̹t�9�Y`�<"�?v��0c66����?!��#9�f�W~,J���M����"���[A�'M5"������X�yP�7�������|üY��Ӌ��������SDߵ{�O�s)1�L����`�:t�&�B>�w��_���4�4~d5pDL5��`U����3���A``�����y�m�1��'�ǳ�_/i3tdY|���E��1������h��{:������1ں��Z��t�飩�����ա9z��q[����;|d9f#�*�' �2�bJT8�UbۗE2��-^E�pX=wR���.*�x#��6��i����gZ+2O��X�曻��xN���pG��n9ͼ�G~�բe�~�(5V 7#���o�-� .��ߡ39���q@i{��|�O�&䭘5ɔM�8�y(W�Vf�5�[�⾁�}��P��k�W+au��3SU=���I��?qCݦfe�1���a�9���4-�c�M�Z�Z ��-�l)�c���r�/M�FV?�%%�ۧ�Qt|�
��W�a�5k��Js�_��O�c�]�2�y_��ؒ�\d�5���)>�ء����9z��1։�T�b�7���A�*��F��N#J1E�m&A7!��tl�}�D'Ꜫqӏ�`�
6�Q��:`>?Py��TEx���Ny���)������El�x3������>�Í�����DiWQ����s�Fo� '04d�rL2r$��{�M��ɶ���*�w����%D�2���&�萶N�4�����*K`ĺ�.�.3��L���i����k���nx�%�K��r̗�'��(l >7��Ї5W������x�{`�>��;%�U2�^0�`[h�J�*�2Թ��2Q�E�|3�uIN��9��7Oc}2q�0�D�Ww�p?:�!�eE�����G��9@�n��y!�I��'gt_KFk̰�&f��(ȫ�/Rޠx^ ��Y`Pl? .���p��^5�z���Z���Bac���19�n5�p�����I�%�LR� ��40���r����Q� ��
0�E��u��VE�h�M�J��t�e��L�i�-"~ ɂ���=M����ޮt�����-BN�Bp�������d�Ѧ?���߰�9�b	����J��PxJB��9#�����0�fڥ���;�"T�|�RV,U%��^��@�oI[7g�.J��C�u�+<���6���T��X�Zn�]�M Jf����M�N���Q�6��ؔUAU�<Z�� ����|�_�W�2�^�Y��[y5�����2��JG�F���߿NZЊձ
�B�?,�H���RI	�u���9���SP栉��aQ�<�Y�R���U�t�R�L)��H/d���x���p��۵�����*G�`�;�����G�M�/U��1H��)�.*V`7���i��������.ln��Y�qO�"t��n��?�������4!�R- eJc���	i�އ<�(����^�4�p�!�[&:}�G�z��cp�4MLY_VQ�ŭ�M{7��}~W1�lt���������. ��=�Wƨ�Q��<�, ��h��k��Y�!� �\z�"�&v�r<e[q��&J?V0�ܶY�������]&���L�E��E��O���t��:�jL�g���]�5/����O�XA����;H�e�����U���_n:�!ݜ����4�#��;�	���M�lRT���kڣ�����4:{?֓����\�@� NK�q��n�zI^TQbRWgz��^e�~n����=�E�������!D�9�1�ƨ#Nw�I�ZB(>�������ߧ][\Z�u��;�s�\��z��o2r��	�[��������;�����kBD>����!�gx
&A�UC�_9`4�ON���(0�
eh+�l%'�U5/Qz��8*�l����&o�A��rs�^(װH��p�����4�èW�΢_��1�����o�Pb�~P�����0BWo��B����:���l~�D��`|"�xֵ�G��z���Qq�"���/��>� H�ӈ�e:>�ـmI�bQ�a�nZ$���kxF���B�S.�GO�s�2�ְ��f�@�1CǊ�D�a���+%D޿Q@76�6�ƅc���=�vo�q�[��&~���%/����}�و���x�!X��#��8P��Sڦڜ
��Ʃ�}��E�I�n�,�5l�l��.��꼞/Md4�}�vj-ҋ�����
z���a�fnrm�B�˼[�Ǟ����jTr�. �|"xen�6���NOQ��[
\�����6��z�Qd�!D��m��΄�j)��j,���q:��G46��Y�/&��3�
=�T�{�E�fc��\©��Ө��O��S�R$ǃ{�K��-7�C��%�h����<C���i�2{�:���
0��l����������t�
�����6~��b2N���C����+������"[�W���F��K5�9�_���L)$<�!�hAS��V_���"�2��_[S���v��7l�����k��c�#�:o���p&W��n�I,K}a�<�G�Xs:�%�9M;VߋM���qc"J`�ر�>�4m��>�-8I���T�!��L��������DTAS+��Bf���xF�������p��ڏgd�l}Y�p���N^������TSjwn�Z�`����sL��"� �����LKAt�9��(E_Ŝ,��8�J��=�wYt�W{b�2Ӟ���0%������n�ּ/�����H�XkL�a�Չ�Q�"�äw`
�f#�`ZE�x�R�	�����R����q�p� �<���v�!$����s���lh+�;Np�~�q>M�(WL��̥���PG���Y�"��:�t��CҮ��|Џ����넘7�e5h@�ڊf�DY�,H��,�cN$��$]���`�&�T"��u4."��{0��W��\ԓ0#�X�jA/�$p�KNrG�;9��չP�E`���p|����<�>7�_8��^��M>;W&ٳ�@��2L��	D��3�����H�$�U\U�O3���oMڈV�t�y_XP��Gm�[�����������gԜ�����Gq�Ax9��-<K���Z�B�s�a.Κ�SD9��]X��>B���
�������np�T�:��ޝukv^Vـ9�C6o�B���N��
���)��+��Vߨ~�����5�c�5�v���'t$�{��F��־�W�ɇ
�2B��Z�p�r|�3(���qc����k�n;�Հ�u�pk������3�S1����]���g+ ��W�����w�x{�i��!A�L{�!��n�(��.�}6c��L*��wH�/b9ո��%��F9e@oI�RV3~qD�Q��ͭrT@$bc��a�����8?�Xy��="�¨l�%Ƈ��|TE� "�P�?�_l�^��]���mm���c�x�T�'0����1�K#%>d���82�2�.o�}�_!�L4�p��4y��-*�D~0EHi��=��/IM#@'��|>��]X��D̃Db�L����7^ý���ԴA��NMm��}��g�~
*���#����+���p�r�N�Xm�郵��~�n}ȵ���aС(��1�aq�p�Bo�6�����Z5�9��Lf捫�.\XO��{5�"ٓ�����1cVL.Gr�E�0��\���Z�ˎ���J0'F�"��%(��o��3���H��nK8�(p�0ٹdd`r�42$#�|;�K��2�0h�Ў��[�`�X��C|�ܿ���D�Z� ���}3�1��.����r5��"�t����и�C�U!̢�����9��X��t�Z�ͅ��K��f3`E�sɄc������5�DQ�1h���pp��d/fU^@�y8M-��`]�]x��������sO���NAǠ����I����A�Z���7�����Do,�����/�]ac��g�1��������ݦ�y��ȕ�%�e��=�m4̄�'zKWd���қ����
��I�{��HJF���IE�����I�RZ,���/�"N� �_��02����p�'����!�5s���\��6]��D>\jɀ���Th'����G�v&4�l���bǽݾ�MՊJ�[�p����Q[� ��ح)�� uA��C�����­�^?��X�=��B�11SΚ�@�,Bbu%!��LCJӥ�զ��B����#e�rmQ����2CzƘ��Z|ĕ�Y���~�����Ņg�d�`�K�O�5�bb�sKm��w��+�O|̉NH��ǩ �d�NUzpe�[۽�]{&��sr�R�T
%
y�4��У�lEf�vu�;����(�iG�;��G0׍H�y���yM?��WH����hO�-�t�]ﾭSI�lN���V��1jR۵B��4	׮3@��,��R�2�Q�'��q�z��(꼋G�m�ںyG�Y�e�Ep/��1�b���(��XK/��_�{A�p��<��l�����&K��R	�[�0�^]�jh��n^RZ_�	J�*G�6�Ԭ{�b����gK}ř>�n�N��ㅐ�kV0kV����:�8�%��˪����k��J���Z2�r�9=<;
}��*J]�U� �D:�ٴ���m�i[���hˡ���[�-��-�w׽��
B�a����*��1�0DX��5���jwHF���q��%0js���U9��,�p>�R�ϒ0��O�ԋ���G�&�c���F�oT�^��y���B��0q�)Q�E���x���
d�&k3��B�����l��=�h���,[ �Y�H�j�˪7:�iCW[��v���`N��x�2�_8��;pO���#/m��(����`���H���*�wð<��~U)w�3��)M�Y���m��z��٫B���q�����40�G��Y�f�����?�)<aPCY��5�]'�k����}���-@3άf�!a!sQ@�׃#I��A�:���%�w8�a��~k������
|�����H�Sd9������7�����H���h�s�Zʋ�{���_�e�"�w�n7�2���҆R���ǥ�����s.�p�N��a�`���X�������W�1zkB���=�����q�[�O�>>��a!�@h���d�e�nkL�V2�`�C7�T��؇
�n�i�\���0�.�a�kv���:@�:���b��tF�˭�tD��-�{w*C|]��B�Ƞ��i�U��'�5��7�:�I��Tc�I��|�a������`���p>M?�P�#�&�E%\�)p}:Va���w�7�Pcv�*�E�e���W8~�VIN���ű�\�'��0���+�Fט�TcF�r�݃��4��q��@ݿ�d���(sØdR[�7])Ciᘡ��_��]�����#���57-���I{<�"���r��Ȼ�o����8*kx]�M{�<�C�j��v�ՕH���P�*:{��� �U���~Kd �d��y��\flR� .R��1����ң#�ñ�����m���1_�g����$���
+�'B!�^{�3?�c�'�]��J9�=f���X�2my�	E7�x�g$�7��Ş��5���¯$u�N�3�jax�_��á������β�:�;����9-�(��1��8MλR�4�C��.�1�z���J�S:)Fv�9�i�Ro_���y�.�u'�t�:��e���~�hA�%̪յ(�7��n8�B���Ŝ<������xD>
/�Ou��!�Φx��;���
���l��97��SXp���)��L�^�V���9�~��y��@�-�&�����;�3?I�Db��Z΃"#��0�*��C=
���S��
�fd8��1iQ^������d��������T/z!6{�V8Ovc�$,O�e��}��{c�r�����]C������u�ꏟu�+k�m����G����|��w�c�xqRL�mN�wl�1I��]�J���)*�����g�ԛ+�J���'�aQc�9�=/�΋2���u&Y�����~�FYj���_�ݢR�ڨ|L�*�f�I½s�
G�{ٹd�>Z��(���%�_(4{���M=��~��}A-ўo����lǅR{�7���J'�[�>��ᓧ��hy�D@B�5��/F�*ͧ�^���|�A�����^9�<-L¡� V�H'*��g_8���4eZ[��ޅ���0�rΥ��
mG;XΕ�c��u�|��%&��ࢼof�iר�n�C�<�rs[� վ{QXcП����qFh�5�씎�,�V�N���zC�J����U� |�F����J<?6$��z�a���<L~�T��꥛DK�D�r�n���`�����&�dP���}�W ]����H�z}b|||sJ|��}4�E�+A�h��6��Q��|�WV|����uz�ͪ�6K2��o��m�Oll���qpM�N�-��2N�WNg;���o�֝D|á�]!6Hΐo����T���Ƙ?�-���班۪G�$�y��y�w:_t��؎l�2!y�z^ͺ`�x�n3��^��0m�җ�L����5�����̬��+(�  !bC���?'��ˬՖ@w?Kj��cHD�_�-Yn4=~��厚n��!�Z�d�ѿ��[�:"e	Y�>5��v�X��t^زx����B��\�Z�BUP�?8�1՝��K}��9�g�N���-����;b첞���X@���o��/U��l��߲�y51�q]+K�.:�c۠��F��f|�i���C��a&G6��������$�y&X�v�v
"���g�3Kz@{���+V�E�]�������7�۴@ۯ��!���:y�z�%P%(%�ǈn��Tg�T�l�p&I0F+�
TH���h7ޓ��Dm��PyeyT_�����3����pD�Z�$PT$s��5F�}�Q�E8����km�0t Ưn��"��=���؉�x�e�X�Z��b4��k�NEw���!lz蚁-��ɮ<Z�N��@�g������$?���_q�����,�/�#C����-=g�۝7�r�?������P;�%���X,L�n�������C�g^z����l�X7�l{��Go�Q�z(�G��[�a���[v���^(h�C�]�V���g�t�����48ꁾ�P�����7Q<��r@�����$�Q3����8��V<�,AX�F�[{ :��h��m�����r��ݙ�^��˩?�x��&�4��j�.��ᡒ��xF���Lx#1\��ډ4lT�c�����Ǡ�d37�,�M�����'-Ͼĕ��e��yy�6���^�$����3�i#{��L�H��w�^�B�bG$�f��!Rfߤ�|SS��y�,�3-ZD�F���4É�D\PIڻ�g�Mg��$���a˼m�KG��~�pL�>�k��K}-c�g����Nj�n!X`#���s~��V\�g%�]�&f���rh+����t�pZg��&��M^��j���7�l��ť�'Ǳq��?�Em�w4��L�\�����䥗t�8�S8���%L�O��f�]i����y�3V�`7��/B���n=O C��hvJ��c�&��w��GVx*��?�s�ܹ���ĩ�ܥ�f�/>-�'-�|D��^S�u�1KB� �tH�Y��W�=��"�Q�2T�sڈۃ�>(Y.Tz��>��A6��Q�re맃#BҨeM.�u��5_FA�_i�ɭ?�æ+�ˀc'��,b�YW�?F��0ܱY}:�����_���7?�J�Aux���,G����ҙ��L��&�}��s˭Ȕ@ig���(Ȝ���!?������,�Y�=����;�8�(�t�qw�����If�B�!�Ь|(�@�&�J	���Ia�Y��!�&�ʝ����ԺX���i�|�>�P5FD��
�;e4l�i)��+'���� ��8����Պ$@s*�#�?�ƈ�4��1r[�Ӂ�9�}7��(v�V�R�Q��k�|�Tؓ��r�g�3*_ޒ���KS��Y����c�^�m[j��I�+���E{잾o�����=y�����@2�P�=F�`�S�Y��#��͵5��K��f%�	�Nr|T��*�F���\&C�RQ<�@g9O�o�3�Q�͛�v��,�o3��-o�9���F��P	�l���� �:�@�E@�7����������qx_VR@W��=sWo�����J�7�M+�;u;)��S=CN��G�9�e��ёa���W�=<��j���\=���O�H�W�"����_�b�Ԓe�0L�Qc��<�O0D�]:v�gG�J��+XPk, e�ޛ��[v�_CF4BT6Fx�8�&f��ms���ә�T��M#¶��ٕ'm�J-c�T	D毋�҇�wr	K���L�W�
�q'�����*@���*��d���w��ٌ} V
p��_@������ч|T#X�N
�+g�����͋�}�)}8��ĨFCjS�Mc�ʻk�OG��/�F�o^�5��\x�Z�fb7m��	C���B�4��	ɀ��^c)--U'yј�����A�J���� w��S=57�� b����%E+e��}��@���GdE��������C ��XC�g�u���û}!�ҟ`��S�������n �9ό��X�O��H�fk�A����>D/rf�lQ�S*������J�FxA�M�2���r��j 2��e�5CO�������hv�*�6�T�s���a'�5{ ����kROez��*��ԋJIVG�"g6(FO�QF ����tjJ��)�x�����V3��xZb����5�a�f(����T���}��&n�wK�(A���$`�) �1�Wd��������Z���!�3����7^��O�&q���OKn���J,�8�v�8��UR����T���fϢI��ށ�/T�
�#5 �N6�D��v��#�� Њ�������a)<�gN�>79����
Ȣ>�Ox#&���d���p�`������NV�K�KN���3��\����±��va�}����g���� �k�`�j'�����<��<@͒����H�#��S�	�lqr��Q.n_�}A�B$���!�3
��/���W7��OH��R�Ach�p��\)KjT��a2e��랲�G0g	�����	���61ۻl�ro��b�'��⹡��� ��^'2�G���jT��y�Z���͒0��ow�=�skSS�P��=9��mJ��UE9�hۧ,���xDHdK�~�Q�N�p߆ l�&F+[�}�V��ȓ�1~�2-Dbbqa�Bß�H��Ӟ�]SG��˱x7A����WE�Zw����f�JA��@iH��	����"�:���G��=���]�=��O#���EGp��H�P⛲�Ba63I�f��d���t�%p�����"B}io�����c\����@7������ܐ������U�������/�oێ���i�n�<3��F�ޤ��%L�{m��~׸�֣��QHw��?K!*�f'aC.UFb��즫��y��Zp��:����
pnTE��v���s�����y��N�S [�$'����M;�Y{)E}�GWٴD�nlsX>AGSb� d�&�Mˇ�OX�ٲ̊��B�Fa}����{�?�+д���#$����tƦdNޣ3)�b��G��Ѧ�>�:�㾘������0o!d����N�Ya����(rl�%��(�aW�KPUR�ǴfO! z`~h=�A�����%��^ڀ}���;��I1>������]A��>��G��I�m@�iF�\�7�K����E�Ũ���|��益�$_=��ѐ����E����7��M��6�d��ma��5��)���%Ǜ ��T��y��h�R�3[�A���6���:㈨��b	(�ٴ0T�t��[$�*d<S�^9�Iњ)�+�3:wؗPN#;+�L��=H�V6���@�V�/ą�&����.;�����{6��)�c)˙�銀0��>5Gc�b)���B��0+
�Qk�!GU/���w\�����U?�nFv��K��[60m;iV��4A4�b91�3:��I�t{��Y�&���X�qzW����#y͆�T�-�#�F	&*���*��e_�a�5?H��Xj�:��h�z�� ��I���b�tVG��S�3}J��_i����R{��"�#�S@�3@F�q:'|��l�O�:�'�`/��7�e�D�s��8���f�Ir� r�K^�曠[6�U8s�J�S�b�'Н?��Z����� 2��BIޝG�pFV��� ���G�u���2��n�ה�s,�,RNuw�)��Qy}����u{�Uh���b�ڇx�}c��m�a��HV�Ah*���e�=�&vFl"���c��j��Cq8��������faС
J� ?�iJU>��D�a�/6�f$�����2n&�(o�/5�
�)�0=%����M�"�{Gj���V�4)k����#�m�@�� F��a�`Y��8z�|�k�b��������o��<�g�&j���ԄcD��qp[-F��؟*d }�X�.�S�5��}��\פmh�1cWw�#w,��{آ>w���Kg᳷�w+���0�C�
y��Bp!�`d��=A��,}�5Dڹ0Lh��5R]I�j��m�8�� )��U��d�����\�?�)ޕ�T0C'ܽ��H�bĵ]��U?P#�~�,��h��h���q�(	ƃ;]� �� }i���J�.��o�[�p��-��+���)Ud�3���_eG� }yW~IŒ^J��G#�}%g�B�G�-�����?���';�fZ+�tl��ԍN�L��)�P�2d�Q�p�Ԍg!Kg���YPe�u��_�`]��7�b�mѱ�mL�麝�V3`�(�&�ݱZv��	� 9�������2u�l�3-��Cd�h�k��opOM�Bz	��R�Fxz���L�t�/�'Vx��K�d��:�C��k�H�oKf��yWf�B��:���l��7{��̧���zYW���CG�z`+Q]T����7�M.K�ُc�vK7"g9��Gpج�����ؐ��v��������%]M�x�!,gy\ۅo9G�ʬ��c�42RBPv�5��*�ȏYr�Π=	�֝7��'�4�W�Ԅi��r����7GG���;�itϞ����g@���j[в`���"Z܉ifQ����g�����$��