��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga��ʊ�tl	]'@q��������M �F��@H���B��8k3{�B>�1̧�^u��%J����g�J�zh��J������	�U:�x�4�C,8��Ou�b��J�NUʹ�vi�Q��3R��� �T��MpE�X��g��	�,��Ga@�\�����"kh'\��u����������Ypqo�ӯ�A�R%��0Z�ƴb(1Y3aCF�@:�j�D��i*���
������n�
�%����w�%��O�� <��k9n��%���e����J�U\��3�.ϗ&gYw��f������3y��v��N��Hۙ�M�H����T��ą�8�9��P7���l�c��,��,ɔ݇��tu���%~{r�le�;��2�i)�P�}n�VG+��-\��M�RY���T�*b,+���p�|��+�.��]ȸ;q����ʞ�\���k͚��
l'�|��a-�٢�飵��<R��֞�Z&imRn����ҡ�����!�����ki�V���/�-�I�l�]\�龡CU�@��H�N�Ԋ�����E6�gD���5��1=��v Xj�m���������/_�?�e�<���4=?2���n�ʭ�}z蹾n�hpedl����A�����ʢ�S�yK��zz?|���D��wn)���o��Q��� �����S����j�1O�0���U���u^��v9@�#H?��H�1�n]�	�YL���sYC����H�֭&7������\GD>_����ku����9eo:<b�}jw�Җ]_bT2F�����Ѯ�E�~R)�T������ v�e���y�a�tg|燧��'��&-�|BQ�AEQ�l�Y_��%�E�hk��2�~ˡ�ZE�t��J˟P��u�ݝ��{�<�_$�)ղ��20���K�����=2���ڞ����ޡ��4<�Q`q�����}�8f�$oQ¬��A�X��B�v�Hm@�]�N��놂ȼ��#�Ȁ���N��^�W��l�F`���m���V�7���q^�%�E�����tXj�9����&���L<s�'T����*Z�SO��`?�a*$�+�N�г����O�(jh�t�<sr�Jh�Ʀ���#���9Wp����Ю3���	����t���[�^
g�?���܅�I�~�n	�c2>�J��0��CZw��5p�>��w�b^���p>���ǧqs�'�}��f��b�6�*�p���N�H�~��DWL�|)��[b~m]0mt^bZ�"��qu�=qqe�-�>@y�9��H2�����(��SE�=��:�uF��K����D���v;M�#?-�DgJ��jGPM��mqW�O�������h&�E���FXCfv���m�.�l��R#Z�7L ��{v=ؔ���w��펭�����Ø�,!f��+��f@�m�9�lqtj1c����֭RN��j�s�Ի����UC	���	&+l`�����" M��KI�\t�jS	�"=�-XJR [��*q��F�M���n5��INyw�Ā~���������j��~;S$U!M��,�������Y#���7��9����*B5h&��jI�UM�%��I=�qW��W��*gl���X��%Y�6Bޭ�Xۀ������ÿO�CKS��@���_�b���1 8�w<�O8�$�j�S���3FQ��H���5��w��:,�ӝ��1$	�-�ѫ
�����	jw`����ٮ�n�]T4�vs:9uB#A��'�i7�e��K�قeh%�.@�h%�yhd\N��S$�%j|U���䣑��XI��ɳ1z5����UC�$�a�'g���.Oa�ʒ��[*�]��)1�������l��LK��CU�U�d�.Q��H;�;ƀ��!�[�(��z"4��Z���z��~������͛��Y�)�^��RʫF����Tk>�@��*"[���$�zQ���-�Dvâ��D�k�p�rH��xx�y�0�h�b�V�{�3��.~���W��u$"瓡i	@
�W����Mn#�*/6����������{��o0Z�d�ߜO+��+v 4�t�Z�	"�j��_��Z���z�S�t*8X�p�U�����RR�!��j�%ϗV���=�精���bWrF��,¹�B2Or(A�>��Ec�r $�Ba���kM-E����i�5���u�s�>D��C$�k��[i$���LZ#��ٯD���(n8�\�W��'����2?U�|6V�Z_���B��
�����pY�n@�[����w#[���{+S��? _П�n�
m��A/;P�I��b����-S�[C�݄NȚ��GB�,����|o��x�Z��A'��Cs�4:p��˾��q�pF����'�IƔ��e>�b@�!7�_-2�)���-e�ڳ
AӌP�sm��������*�Y�:&���^�ohm8�i��~3N���Q<�[W]�ZU#�H���(����DR�*a���S�ߝ�D.���#'==35|�Q��d#L�/�����ccɤe[m�.��Z,��k�oet��g1���`�ܬ�R~�xl[A�C��1�`e�;t������1�:e�c����zOփ.ۋ޷���s��MREp����Mks��}a��l�a�1{H�h7�p�^���^v��Ư���=��m�8k�Qǐ��n5���X=U�ۈa(y�9����.�8��>�&�y��N�&�{Z��f^8��\��k�D��\�yNdhnf7��0h��X!i,�z��oN	�H���P%k��~aro^�,�#Ԥ�B;���R��Oy� �p.mku��m�M�XH�^��ݻg:��%�ԝW�t�(��-n}� �@�QZJ>E��WMݾ};��~0^e~� �}���J����~T��:gYk�	��ə�C�A�����7p�CC��Eo�����ɲ�S_W�����0I���F6B/�	�:$o���:��x0T,i��O�X��M~y%�Ř�̰�K������]8�f��M���n�03�(Ew{-�����Q<�'�;�γ�n>�A��O�:�[���ؚZ��nE���;�(���3��XYcQ�UM�׈~	�`���y�������J��p�u��-������g�&�D��]|eX�an D��
+;�L��>*�r�Lh&�ٕ�'\u��Cs�%#�'+d�7�w�Ȑ�ED\���:d@e�yB����^?��^�����1��F���k��09Fd�-��7-AS��_nXR����c�P"H��`Zo/�l�x����6�#�i�6� f5NBI��:�>BpK��um
-����".g�/�$��Ȋ��D�<�( ʛ�(�Y����B<�����	�w�x�����h�x����V�}�$h:�j�$喆㚥uE�����#��0���Q�"�5�0�J�;���W[�T1�!S��&���6�Ȏ��Z&�VL�R�EH�~[�a�w��~�'�1P�	�{1��H����2�ڙ�څ+����zӯ�iC�έ�PB*�?��(��<�؇�t%]���䙇q\�Z�'$�1o:i�#�56������7����\��}L���Z�i�>��tѐ"�W�B��86��9�bg=������&o(��&�^r��T�QX�����`(P������=�w��w>[��XFr;H�������ov�/_q!>�bn?����70������?hL�#ǥ�ijU
���^�a�^�g����h����i��u�� g��ԓ5�y���䞬��SWBj�~S�Z�JHsG���O�4C���S7/h$S�⼮��	��-]S>�bt(��	�*����|�
wZĹ�9.P�*�ʧp�_��=g�n��ϧ`oˎ����a��[���{��W��R�.b�+��п��;�� >.��&D�8XX���v�~]�J��e��86!`��n$S-��;��9P��Y����
ǉ3l�R"8h�>�����T^|����!�K3���q`�)�Y��j�ր"9�ޤR/�k+�iU e`lȻ���+���(j�v�RJ��a���D� 9�X���@�a�Nb=iI��+O�h"�L�����O�7n�ӔQ5�(��I|@=�W�c+6_(n�p���	� /��8i��I��:;%
� �|��:)�
DGѤ4A˄��r;��x�R�y]u����1G3�9�p����bБv�<f��,~#��Թ��"BJ�&�H࠹�¯8����] EJ_�^r �r��=�]��R�fg5�"���/��Y��D�������Z�gt)�����Qqw�!ق��U5t�r ��'���|m�q� �:'�@�T��+�͗ �J��#�Ɣq���q�!BE��[A������e߭u]��A-�Gz� #����(���i%���ؖ6��s�����_ȵ����D5\���OI_�wy���p�n��1��s��0��[hi`��1M�q?4��{K�e�l��	]�4�a�+K��ϽO�Yr�R\VKw��^�b +}�lZ���߉����	��4s�����:C��8c{A���q�D�!��OϮ�3��w�?�;y���R~�;3_`�����������ׁ���(ATj�2m(ru��V��������FZ�7�;���TQ3����Y���Ó�"����+�����7+=�A�����9oA�4D\��&){vM\O\�q1�T5�.��Ϙ�`s�Sx`�%0G�n�_��Y8��I
�&x�R,��MG�
��S 9�?�o�]�r�s
s?M���t/�� M�qrMX\Kj���zw?��{����m���S�K���x��.�󳩎b}4�ʸ�?�ƛ�36���Y���0m K�Τ�]������+��]�J^��Н0�5��l0{��Ҫ��]����6�uDLRb�uC����k����	�����\ۜ��	����h�8�v
���OJ�2�-������o?Hhv0�9]�eã�$�h#h���0��&<�C	�9���[�(s�cE�쳯vſ������`k�k[BY�[����:JX�_���w��5�N�y\�	���ɑ	?&�����bǎ������b^?��Q��]��i'��[��߶��2\��#��8�q7�];���t7�U���pGL�m�	J|=Z�cm���C*G=o�+��8�+漶�&� 0>��S/}f�����p+��W��~�E�}� l:�J�����i��9q�oᯄ��Ƥ�ݑ;�-p����R%�nu1m����*�b��I�{DONs�۷=�H5�����zѦH����U��Ӄj�+����o��^kEn}�UF-|�dçl£�H���N�����X����Zշ;���0�Ho����!fo�m��KU��֮NN��U�uz���Y �ˍ ����r֪�=��\2�Wtꫤye9	ۼ����Y�;���3i�i���jl�z����'g9=x�SF?�A�*�/����4�0)�V(��(+3���V׆��,��e�ԓ�C��(����dVױKJ���-$�!}I?ơJ��wL6*nq:\7�H�w�C�{��}�=�b��8�%�]�����9��΀�o��S�]$x���lD��[�c��y}����82���4�NC*4�|����2|vr�;,L��]�<�!�lbխ�)7���M017Q|g_�Co^�Az������n��PՐ����7"`->�O&uD[/��`4!�l@�������F��G��[2ҡ�����M�w���gvE��yop\>ǚ��k�JSk�s�ٖ���_X̭�p���6ɐ�(�a g�Y�͡8��Ǒa�z��(F_,Pm��>2�3EcA�9C�#l��îe|�TE@�:���lD������~�6��OB����]�T��`�r�:K��!�Z���F�%����шS7�&+�gX��{�4=s����:����{}�{�]�u��
�����͝�����cL'�.B3?$z�v�Y��3�Х���a_�B}.��`x"��A?�z]Vm��w��;��3Gwᕣ Q�be��ʯ>	����%p�{�[��jq���_u��!��F��.�0� 0�ҙ%!����������������D�Ь_j�H�r#��e�G����M��yNOė���*�t�M����a�yTv��3о�&\�9.��������尔4������eJ�B���ӝ����vo��H�vN��Iu/���^Ə���l4�ĨW/��^@s��w����̖Y���8�a��9���ȉ��R�����C���-c���-L�Ӧ����:�'Y�l8�u�.T�����c]�י���W A�s�eH�q,$����M��1+vN����K��ik�n����� �]n(o�Հs�V�u*<Yi��6�9�P`�f��ex�X���y�-s�o} `&�V���A)bM����P��(�{ҭU�h�b�"ޮ0���1N[�X�
+�t���Y��0�}4��=��k�N%�Ć�x�BZw�ʼ�r��>@��2	F�����E��L�
Z��3ZG1��b֧��Z>|1ѧ驊t6�
�ÿ7)c�C	h��q�QNq�7�<�DH���	�x�&Ω���Ω�#0�W.��RZF��ۋ��x�J�Hc�,��qi�n�|yB���w@�JEI��9i�����,&�b���3�k��^H����Y׷ȓnt�R �?X����gz={	�Z
��g%U�G��yNtɶ9D4|��|�_�`�eb�g�����5�K�g��qf��M��K�
�V���0��Ӗs��G)+�ЙL���m�hN��Я��I�)��[@j���܇"�nP"#�b�s@���;P��w0B����PN:���o��x[evF �Ȁ'� ��S3^&�-,�7r�v��a?eZ��nq���o�!�w�q��L���Q�]m��ށ���P�r���Z	��B�f�~�ْL�����=v�'�J��-������o}�h�|���\9ߜ�=Zp
��auP1L� �)��dV�VN8���(υ%z�G�7��:a��)��G\�h�%a��4ջmwf�
Q����Z���(�|գ7�f Y�c�;@qz�>Y=@{my��q�81-��E�^�+8��2��r<)�ж!�������J�$}E�ty�O��H�s��m8_�U3�uc��3A(G>[�z�\zI� Z쒳���$�Zz���/��|��� ;,jdd85��_����%z�?N���W�k2:D8�4���\F�@h�f�W�a�F�6�|��@��)��]���̸�Aj��2j2����_<�I����e�G�|jl��MҠ���0�ݯ�1�aT�t��n�);��r�}��f�Y�����������%���i�����S����
CB�:���T����z�ҟ�+��Í�}��5xQ��.j��r�1z/c���#� �ey���O�ʐɮb����?� ŖBQ(0��j	"���vx<��g�$a�7|�ڽ۝L��C�Ɂ�o/��n���#�j�4��kN�zǤ�R���'ac���:����Ҽ�ۃ%�8�Cע�O�ĝ��~&&��FU�8�_l�u�f&!v��wH�QP�S�r��ym�V�'��>J��o���t	����6���ܤ����w�		�;3�F�$�覎�Ε(
Jm�/c/���.�2�=�C�Y;H�Qd�.�x�v_j$�9�n�0�MA��Q=�t-�����lo��K.с!�x���&������,6�G��)R��+�?%�3��qr���_�����K�t)�mѢ�W�F����BҨ������jz�'��?�ϭb�I����WY�/�SL�|hH���-"(˲��,�IsJ�dq�!��j�fV_R��a*�ה�[��ϙ�
w�G;�'��@kz�i	*��֛��e�
g+й� �bc5'I���8�ĸ�YR{Y��h
����O/>L����� e^y�uE��?�n�K�����vl��IA �RR�r��Rng�{TWH����7���#�o���"�I_�eZ���9	�[A��9�g�� �"7�0Q�oڃ�pȱ9�8���t�<�i%��d�	Mk(:��pƝ�f���A�D|����s�Uu���x��e�0�xM�+E#G/\���������r2�K��!�26Qg�dD|k���1a߯��9��g
�Zu�:�,��L��IC*'��}Q_D��c��}��92�w2�����,Vt��� tt��Z�f�n|f*ϋ��fˏ�s�i�G�w'�x��E�$ع��2UFP,rw�e�y/�_��i�7U�P�6v�)������O҃"?<���|��U%m���N'�܇*';t��}3�xu�
/���B�acܺ� 7��f�X��*T��	�I5�m6U�\bO�G����z�Q��O
��H���aᘳ��RC'�,����$�l(ʢ��	0Y
�æHw�N�#�e�_U��>F=�j���/l]	#c��u�u� =/ȃ�w���/m?��XTx��6�����@��S��_e�(S�%RL4��]o��~��cc��P�~�7i�a������s5�M�v۷�I��.����Ф��`�=4I�Tk���8�[������2X%7�$1��S������NVj�t�R��_��m舰�z����>��cJF��!� ��m�w��b8A`l��L�]�O���2��{������B1�.�ʨ��T:;mR��p�)��S}���ܘ٥��`6�Mp�J�h� �l4�W��i�GEns��qp��^��F�5�����fL�/����)����b��A��Z��/�=�.�O��T���w��J�z��-r��iΧ ���S.4e�M9�@�=�H�p�0����vX�K��s�"e�/�������1}z����3�S�E� C��:�o�ˀ�#�˗��ҩ&%�ќ���M��0q-^�ѵ��4�_vz���Y
,cR����Պ�k�`�w��9�CE�r=�+W� �bBp�{R��j�!d+5���!���3�êiԚ��驨�\O�N!�@��y��Iɖ\�����t/�_�l�Eܾtr��ë����suE���ok�,!�L^O�k5(v��о�&�r�6��?Ӽ�#�kTʪ
oɰq&�*O�LB%�������Sg�;��a��F�[55�l�j#�IГŤ��ztF�78�u�Q��|D+�򈿔V���ro��$K��&QA�%�H�?���m�5zח�[ξ��9{M��_n��	ZV]!��f���h�DQw��l�?�4�%��G�;�C�����K}���kE-�f|� u�syd1��! q���Fki��R���p*a�A��1�"��q~�r���FI�*��Ac|OW�։}�6�T�:��*�$����r.�U�f�8��j5a�M+{�{,��T�f��y��G6��U�2���."��B=�dKE%h�4�_��&�d^�J�X�p���a�Q�~�x_S�ht�U���DZ�Z�`�T�w����@hⶨT�0����Y�Gy(�F}V�q@����TYD�k��%޼��	�*��S�d�W�K��8���Ki&�����јrRՈ��ȕwM���>A�&�m�[�Gu�@7_��Υ ����ڃ
k�y����ۜQ��(g��Oet2�Uq�C����ud�p}*�c��smw��w����M�L�źo��b?4��'��T���5�+kyq��4��Tf �C�����p�=�Хk��J<$�(u^�����l�۹JEn�=�eoq�c!S��O������.��]������q[y!�+��U!����[�S�|��-w9{�C����(#�Ig(�~P����*�D������Ng�/p��"�Bj�J��R�ܬ��7>�O��(�.m�j6�&��s��?�QQ�B6�_���[���v���a���;%���ʜv�i�K�cYʎ��G�K�L���F�$�z��I~�=�އ��g��|]o�[�ڱ�օ������џAK�c(5pD��)�0���"�_K��ȋ��_���$c�`al)��OF��ܻ��[����%Ul�]͌n�܏���5{�������֮90�T��M��_{k\M�����3�!����sqTl�\�cB���;�%�	��uZ�%�5c�e�V�b}\�U��Ю"Pᚾ��\fnwZ~2YG�5����#���3W`��^�2��i#%�Ri�0�*��L�Tn�o6�g���W��w�V�/��'�!DK��1�Kx��$��䴖��V5�$t��_$]�N���n� �&G{O>=���ɟN�Q-$]t<�OPP-�A[�+O,J�,����������ӆ�qD��a+7u�Y���[�]�6�p��xx܅�v�n����w�5	���k,��4O%���g�LpD2j�5"i�]�H��x�~�&�B'�ϓ��<Vm��2����632���ܯ-�!�5�)y�޹��"�g�/�$�s���'Wa����U33C}z[�'~݂{��!#t��	<V�L�`a9���H�O_�(�G�M�u&m���\7��{�zC/��͆���27���(D���0�aGY&#�dжࢅd�=��UC �P�NJDc�Y�o�������Pp�# V����xi��:�����a�K΄�ĳ�ݑ͒�ȼ��ݜ	����&�L�H�-��%Mr}m��P=_!����Szj��_)U��l.�(�/��a�xmO���7^l���+C>΃�AM��M�1�Rf�ڶ��N�BV�t!��ÿ��ғ@<a4B��	��J�9���p+����2ofS�`��a���J�v/J
:W7�x�(2G
4-�Q*��0�YSף��~2�Q,���/"�H�E�/��B,'��C���`�Q�Ox��4 
yo����A�n�=� :�Ry���mP�� ���wȐ�����ᗝ�u�nfXE�Qq��L�=���̀|�3Z	��D4P�n̡�&����%)���T|��L�$� �*�Vt�|k�����k�)�Z�,ܰm�#�V�	L�?m�yoR��2���m?������e��;���#"�)�Ƶ�y���;�Po���NA�񌿭��&."s�F���t��3;3��1�q��Nϸv�~�+�o@����e2�n>��`�<���N�Wcl^��V�o�R�����w�1���ۏ�8�4$�J�E�K JI.�5<�?�=�	~��6���߀�X<-[ÿPex��ө�c��a�4��Zt��
��V�����s[�b�!�{,)C���o���.�e�Լ�К�R��'�L4��C�Pg�Ü�)��KSU��%�Un�3�@ɝ�uҁ#TV0���� ��{�R��W��p�w�k0d��D�'  |�{�������� 3>0x���ѓ]���`~:�QE۵�yy�s��
J�Y��L�K�5��15Y���QdꄇL*aǗ�,v�f�	Xغ��%�I�
0���w%�[*�� !�s5����"�����|�@[�ʿ=}�5�HΘ���w�s�,z!�p����L��$v�Hn6��o96}Q��G}��t�T5�M"1S��h��н�"m��g��$w̶��w*]oF��7�ʑ��.s���<XOW��*v�-����3�4���D%�^�B�\{2����,��L��{�p�+��(�[l~G%P�
0x]�&�	�|����宲��γlD�ia�P��2VP��τ�ƥ���L�`-1�θhC�,F��p��9�V�>�$�"���X�4����;J8æ,'�M��]��Lq���Q�P1�&��^X+��'�͂u��Xak�IĨ�����C��z��`M?�vAÉ �+D�b]s|�r�4,��E�����'���X�z>?q�����=�"*��*m���P��QY���sl�9~�/�0k��I�����Z|����\����}���n�b��(�Ι'HV�"�N'��kI���c� 
՘R2;��D�?y��%�$&4��%�вb�=4����`�b��ޤ��ѣ%n�kh��#\�yXUe)�0�����!�����(���DK�V�1'�
f����k�x�`���t�q�}�����_{=���� �7��dֻ�l8PA{v�;њ{��ly(Ĳc�}�&a����X) 2��)���O��q~m8F>����ο �����J5�gE��(�X�a�V!��n[��()�� |���_�\/��2uT�J�3ܤ�su���l�T��4<x!(�ʗ>���v@G�>H!)va�4�s���@���8 ���pQ�r�&��_���.�|sk���=�#���'�
���p �?���#��9B@��K���<s��J�ĭV�{b���4��������<�(��"'�Lql�:��J�WC˟Ny��S��j�V�,%Av@f&Gl���V�P���)�e��(c�J�t����">�U��f��f��A�`f���������� ��*�V��}�u�\�KM��Pr=`���>�긳l���ٝ��S�P���L9��A��'i0�o8�5��X�
)��̜��xh�_���5����	uЕ4��f��_�L��Ra�_�]��m�է�����q�w7[q�oa��5Qk��1��s���y�m���U�[)��_������$�,�xh$�u]-H;����}9&|=X�HJ��Iz����"i�f�wb�R���%o�W@��e�ˁ�A��XZ����r�1�N�_�����l'T��z��ڭ�)�)$\
�FY�zh�R�oh�����)9ze�����2Ls=��M5�:2qs�V|�g*2��9������ܧ�N-tϛ4�k�}�u���q&w�ͤs��z�R���{\��=BAHt;{^�rݲ0�\�Q V�DL)M/���&��w�v%�6$]�7V�;d/��rmM���EE .~�e�V�ӧ1�d����n_��:L�\�$��̲��t�w��nI1C�)�B/�����i��T+��!��PL�:Ae�g��Rgr�L�df]�0��Ez]Όk>k�)E��i�x�;��-<���|��ñ����IPD�V����W )VC��PS@�����������k߫������s�V�����+6
���٩\];&=�3�ԥcf�8l��z��mQ%9���^A�B�"*��%��VB�K�uwV�N��u�/�=V��C�D��\�u/(�z���ֈ�p�����Q��ˈH�n1��h��o�eVRa� ��y'�i�»F�e����)id/����J��E���T���D/gF4�@m�J���0XU"LG��|�r�<Ɠ8-߶¤ɪ%��|$RI�3	�׬�aPRc��>��]��JtP��63�f�U�o*��H�P�yTO�5o�J�"I�T
.��=iC&��Z���^�wǶB3�kmsO��8$�;��ڀ�BVmq�,rƕ�y�.H|ڷ���@A�K�e�6�jl{��I���7D�^�?V�U���d���s5���|U�����G0k`���(�+�%��.��ZL
�q�"cw�XP�����Wj�����u����`R*��I�Owf� Ҙ�?� �3-Zq�>����6�s����7�R�R��)
9�?���1�!�t��ڒ�c�is��:�G�E��'���j��m!�Up`K�1��X"o��M]�/z=f���¡���;���Sȡ�w.���,ꤑW����C��2Ŧ��U��&�zX�R���]���z�I�%�����Q�GN�H�$����aIot��{2���S��Cq�0q�K_��D -Br��c�Ӊ�~z©�T#cw�x�X"��f�F؆���cˋdH�}��K植���i������^9�җ�@�o,��tU�
S�J� J$�w��� ��P�p� �e�0��"����+�P1~S�F�r�	1�dJ��&_8��E_��A�+Ӊ�U�2Q����G���F����L���5����E9����E��Sf�Wd�8<嵏7]�A3���39�B��эOt��f�B��IFx ���f�dq=ݲihU�l����Ə�n���k^U�_�(b��"�Ɗ���q��s����F����H���ެyxP9>@���n���&X�Ou��`x>ey_��.ٍ)v��P���*'qI_�QnoSf#hH���$^3�s#�)X��r|�)Eͭ�ǛQ��\���ov
R��;�˅��H?�D���|�u�<j�����X���t��RŹ?�$�O�3jG��e��������#�Zr��]�FH�$Z��[;�S���4M�ח��<3Z6��_ qc�H�J�n�^;E�jD ���n|��6h�Fp�a�Q�p4,�GV���l�
�P,D�½�҆�*=��X�O�)u�_��:�f1)����r�����+yGg�����ݯ� ��� ���p0��3��C���$d��@\]+�O�#ε;��w�Ҳ���N;� ���q0�n3b=s8�Ym�W��B���%�.֭��A5�������Mƾ�
���7�= �їbq�=	�:d�+���*��,0��3B�)�i�D.(!x�e����끗;��^LM�v�$%���A�)�q?�/���X�E?YL�Cɋ���6�ۙLi�Aa����U7J�w���h$D�Q�8��ܘ�ZdUa�lQ��eAN||s�L"�V�Po�$��l���3�����q-(�]�4|�$�*ޤ�7��6_%������c�8E��9i�A�[;/����g�\��$���ư���m��4��6BI���v.�[=ƃqh���3*�r���M�G��{�#,H]�XB���'�9�K��d�|��u��9�bYC���I�)���~�����b�+��(��jmF=��R�e�e�`U�84c�=g�yu�w'Ϗ��8G̹�_py&3tQp�>�0@>�?��p ;L�F���ZKBV)�>Q�[�l@tA6Zgn]��Ŕ��@r[���ؽ'�|&� B�P��_��MiJ�|gs6ێ�;�w��?n�a��G�+=~D�e��E��(�an
�O6
k�
D�XJ���z�\�R	�W�28T���/�|� h��T!.3�X���PY1�Kخ�K}T<���r��
�W|t�Um���j�  �S_����x6���?���K�|�����(6Brz�3���_�O�BY>�����ѱj�T�X
f��ݗ]K��J��^�#0d�m��>�������a��羗���/��h}U:��PMniR0�[��9��PP9��[�y��:UZ�ߋƒ$m1�:���ne4��ʱ�բ~޳�j}}Ю�RN�X�I}`V OZ}�g�Ȟ�,��+��@���`��'��>��d8�6��q�7k���94��0�W���(S^��\�R�K�?�=�������k߬`��(��ja`MZ�jv�!T���}�i��� �{D�P���j�9�$��.i���T(��}CzlI��^͒0[C?�$���&�hG� O��W���zQƎW��C��~?���`�Wc����C�ȩT�G��Y=����"�X��,b�V��R�n�[o����Ԙ�S��ۋc���hR���� 1���{�C� ȶT	v�Ǒ���l{e~wO�N�s!\ M�G�'��3)��¸�]������ �؇S�!��rJ�}������1��Q�_/�`6a��a��'�r�ס��J�?.��7�p�����5�d�ֹU>��F���y,��>	ң6�f��6����	/4��g�;�y�E|v���6�s��ƉP�GI3����؏!?�*KVT�Y��3����j����$�%�˸��A�k�t��Ջ��o3��Wr�@v����x�ԋ�Q�iN���w>9ү*Q�Mq�[*|QJ6D<�O�?nSHU�c��>��;{�R�������=rƠ<9,g|��$�j�DڴSwiI�@$C��������GJ��gma���P�ly�|*!�?)i�}m`�N���v�ր>
"�,�3�{��	�<F�A����:��ز�Lr�}~?�1v�`0�9��S�]k�d�V�e�D?�lŢ-��˯�A�k	�lG����{l�~�P������{�4|g��[������גfQH��	^�d����;�C	-E�}�_����T2J�&V3�����|o�v�h�9'����2�Q[eM�����r��n��?�`h���I2�*;����#��k�"��ΫM</N?Cpe��ƻ87=�ݞ(c�����UvR���hk����4~�t�y�p�	6�*LO�4K��op�G��&G|s�(�t��e#	$&�w�N�<��k}�a��kI�<��$8����Z�K��V�����q��{�s�m�I\�^-��l��[���u6h�ɥ؏�e�b$�Y:`,ն�H�B��8l��!<w�Ƒ~'S{�b��cZ�m��[�p�h�)Ȱ��e���Q4\�/��e�8�~�3�ǎ&x>��V�/vW.*��'�6<��3���Bn	Աۈ+�+e乊إ .�դ�����ۆ�&6�3����7�Hq��O�p�M-��Y��Sl��\?jnR����[��U��Jś��{�]mND<�2"��_w�::E��:� ^Q�D@���&g�_�.����+�_�YG��}�,��3��wS��t0o����y����!޼�%
j�dTs���KDW�.��r C��5Td���O\�Ў�]��A��1|�fTe�oF�D^�� �jG*Q<��m~�jL�.7@��j�r��|h��8AYR�%@N8x*���:��X٥��|`A���3�o�Y��C�����-@�\�K�=j��i�7g��0V�|*5��ĺt��g���P��&̠��qT����7�.�+�7"F�dx+�m�5�V��X�*a��Z4�W��6��@�����&�M�KY`:���zBP�:�%$�Pّ�A�(�π(߻[���R��hG\f�ʓ��a;���=��h2֣�>��ѭ���J���o1���;D5ƭ!���&�eЗ�R�uF	Rh2��9e\�#�%��Z�x��[)_��3�X�9�YT;���֦CF?+S"F�k�F�_�!e���n��>!�Y,wn����� ��H_���i` 4}t�s� CM]��3ۀ�8a�v���ЫIg�2��0O��l�)>UUǊyYj���?���`�rW��u�5n�~��p��<�*��&jwh���Pi�<�g��+���)Q�;�S�K5��8
k�r�i`�,�q��R�kբ6ON��p6�^�-+|ϫG	@�]T�,��W�S\��B����t]{�΀�J�OJ����������>��JDϳ����6��m\�
�ou�.��dSx��t��i���l��.�������_��5㹲�ݧ�a����U"4���q�Dց��d���Eo�Ŷz ��?�~�M:����:���!�q�.=����R��?�"��-��y�`jZW�3Ά� 4�	��ju�s�ʌDm{��t����L_����e�C`i��Ͽ���7�J�����#���i
Z0ِ��� o*��w�~6����!v̰�mۥoI
d5�������4k�ړ}i?E������#�Y &{i5�����%p'�3������#��a߇����b��������m��W��Oz�S/g�K��':�����*3�%Q����}�M�d�<�փk�Dr�d��q��$��7�k�uH���QU��$������m�g����̄!8M+��<u���Wi}m��\xb�Rp�z!�����*Q�D�< w��F�Ϥ�BK��iaJT���c:C���M�)s@(�'/�Ǥ�&�
DY��L��8�c��bL�Y}�:�|;��������"4��vg�{��M5���*ˈ�ۄt����� �Y���Z��##�_P�^!�%�s蚴5�����7���E��pkj����,S�ݠ�/���)^Ϫ�"}��KG$&�D)Ļ� �&t�� k��b���gJ�͊�ݟW�).����M?�u���yh�����;e I����O����]�}���q=b��պG���ɍ���pg%�s^�?V��>Q�J���	z8uM�t��*z]��ud<�:l��5�|X/GV�<N�e�6�����K�i��.b=��cS����Q�liH��B�J��l���h�1�OK���"��Y���Կk�?����8 ����C$!ME*X�w���Zl��N��C��8���ن��B�_7�m�.`.)9�>�&�L{�oε�!������$�f�=��'��{Ad<B�&NHG+��CJE���\q�g^�g��> O)l���棒�	�bg�q��;G	$����?*p1>�yR|�8w�iY��3��]��K�vF���&SS��f����~�rک�����\en_uT���BO�eq�(��E�G#�l�NB�^8�;p���#Ȧ7G�Psho=:�@К� �_}���Z�oEЮ6iϕڐV\�z�!�8����'�. �H��^U�H�h~�-�a��%��
�@�c��&���\����㼼FG�c��)��6�L%d���Qߍ3����E��m�{Ɨ)��"�lw3 �r~�MQ�h��<�9mG�n`�]��3ip�y�/�j�oa:�f!/�����r�g���/������e�y����]嘪��x�nҔ?�  Y��k1p���Z�*W8�&�����E�H�T�Z��g7k�=|��D���F�*/��W��m2
y�Ժ�hB�JV���� ���!�%��g|} s'T���}��,���Z��ih��|cE�#��'��@������h�Y�C�R�!��і��W�O��MT_t5�?�~��zo��@������s�=��+B	����ҁ
gSGYD	��~��������b�ٕ�D��'���W�:ku�m-�	��I̱��0\`2���c-QFҮ�~���`�BR�Z+~Sgstج�!���L�ؽ!A�+���ݤ�!�@���>;�<���h��m==e݇p?��n~���I�&{�(��]�AD7kK"Z��n2�kֹc��J�|����N)�����8�w���V�S1%&���P������'�)x��2�fS�Wk�4��2��[F_Wtj�N
�M0������`������Ѷ�s]�E�!X��z&�FO8���٣
gg�������d�:�S��S���1����E��.j����6�PXF��e�NF.f��g��k׸��΃nzz3<|Vy�m{~Ro&�;,���U5��5���*m�)T�j������=���0T}1���,�4H�� �T���"xX���"e���f='U�dS}���%������5D}���)�n6�N��,����?u��wZAf;�Q�W���R1������lMm���g�+_��>AG������Q������ }���ɧiq��x�I�.*�*��](�l5��Eל�/�$= &��B��.�o��~�e[t�^���eO:���X�0͉_�v$ߐ�C�w#�y����4s"�N�B�gd
Zu���)��dt/QU %��z�3��# 4���<ߡ[ֲ���Z.�Tζ�����eJx����#��H`�k~a/rP�%*r��n����Z�+a6(�[$V��I�j��)�o�C8�����l�IU�)�y(D.�8,͑�Z���_Dup�Md�>�`l�O]²V����[�`X=W���n���Fh�-���
���j��������H8�đ��_���Qݳ�:gZ�~�A3�m�c�լ��C��k���v�X�3�d'׍��ȁ�J
�b`%��d�O>��/תM߲�K���&K��mEZsA�E�}��Dě��{~�{ʜWz'��vރ�fH��U"8�=�tc)��z('	�N�|�q7�t�n�꓁[���f�����{��m���vv�3����)	��^�o��Ǵ݃c�c�@�dTTo�9�C�q�4㓂>��ڿ��զTT������6�Dz&nd�ɩ?����o�Y3�?���:���*�GB-��.���H>h�r�ı��5�ƹ����r���Zk�F��|�K�U�}S��%w�B�C�Fl "�L[&�k�Tk�9�w�oGs;��}�.�Nf.�ɥ �c������Z��V�Lĸͼi7�����ށx�o��{�������Z'�(G��Z���*,�Q�F�ۘƥ2�ڂ��,/�ps܀��n���4��4�*�)W�W$���W���R�|o�;������;�p{EM�Wٷ�O�@�c��K�k�
���<�b�U�I�ڹ���s^Hڛr泆��	�W��9B2��2pu��X��'�A�������.������qX���!��#�����c�@|S��q��+_�Ӣ�Wmʿ%�1DG���*G#0/�m�5�����څtOO��;O����aY$U�7|�p�)�bY���>����U�@Jx��(����F�϶�n�_ō!&+P>T��B�Y��CN��ZH�	5h�#�g�����c�#4�U� ~�3K�&����P���>2��:���S��4��$A"��\�����Լ�kAD�3��J�al���r��I�9J��w0u��$��J��3�P�\W.����|6���Z�m����D���1M6l�bi��Ґ@���_�h}S�9U\�7���F�(O�>riY%3�<�%��Ȕ��͗��,k4�����Hp16%�"��vE�^�!�Ӂ����MI�oF�v��c7z_�!�j��V��}��ƥ'A���cò-dw�Af�+�֤��i��(,1��%�"����^��k���7�e�F�Dz~�8�J[R�5�.�o�u��2|�L���d�m�&��h�)�DEm\>�lQ�Zx���0����QTT��I�"�J�-���DІ[� ���)b{a��6��v���X�!Qߜ��y)33*�BSV�!��	.���ڙ�_��#�O��ʟ��P�ΎB]ކ.o��7����ث�0��=m�<�nI"�eh�	+?n[ssK)!��)�L�(��7bӡisrp^^��.IG׳O�@on���4;N��V�MV���m�@Kh|N���ꛭ�|nN�r�d��5@��+��V�hsn�|C��@�i��;C�O]�$Z2>B�*�A"�� �!�u��vs/" K��8�4#�)��<����o��`�}��w�?cA���e��c\�f<�4"�p]T+�ɸe��79ȼ���J��;pY~��wng�.��3����9O���x��#�@����ց�S'V�:5V���fd�A�����xt��2�0Rl��~���c�g���ŤS��e��1���~���lS��Q���;|�����	D.��s���[����Ŵ��J���Z�=�
}E5fd	r6!�%��ϐL�M
���W͕sw�]�5f�_����v-�|���p7�F�Z�j�����K����P[%�S�A^P��Ռ-W���J|#BKA�c}pB��]a���&t��L�h�-2����h	S��'?���:ˏ�$d~q.%L/_�&����(�[`�c�&]sKn��f��|�)�G���X"B(A랶�2O�gNnot�_?O���3��7����������JG�����f���'i�FS
<f1dQ����a�@��x�½���.������P��Ȼ� JIl�Լ"x��*'հ*|�V����̥鬉<����a"��X��$��$��(28笗�*OԿ�z�A�R�=V��)�Ƕd����27�6$^�8aB�&%�IK�?��6]��5&8NF�M�O���F`"�Z0������Äs����ё��@L@d�9� �"K��ݟ7Jc��5��]&J_�F��@v�ħEa[.��%c��� �0�����P,��i-�����L_�eO����xB�[���`��_�j~��vC��Y�E�aj[$�.�F���*u��_�= ���넿�-K�&}p
X��r����T�ݚ�c`CLYכf��r9��:u4�{B��ڶ1��bA˒^E� B�[-~9*=~2zTqT�
��B��C��$�K��r�E�4H�;��o��mY�?S2���i����*��*6�*�E�p�n����W��3�m���f�>L&$���[�(�ϛ߄gA�]u-�d%X|B�uEd�s�V&�n�J����֮���i�΂�qG����]ގ�l�b�Eǚ�zL{��z}�lε�<�8%�W�H���p�U�����³�mz���č-��{���d3�/�St�^)p$bflY��4�S�9�ba�W�-�/�}�`�S�����f=2�!�?vcc�k���]&��+�1��l��C��?��P�k�C�V� J������������^5��]Ե�XFj��>�����U����>� �:`+G�h ��T�v�������\�Q0A���9�gvye;�0�e@QPii�xw~:�tx�"�ΐ"����x�V��U�u.%JdV��*�p��B//�[�������'R�'��W���+RQ�I��3��D��qls�$�ԑ/��F�c����d2ц�odG�u�q�Z�sA},9K�x�6����_]��Zz��U�Z�����<d�!J3�vx�<<3�������K���"َ�(g�y��ArS� s�Rd:�ڕ"�u�!+*&Z���v�%��x| �e'���mu���:��`���Df��ִH���¨�.���[�4��/ɡ���T�4Af�X:Ry������$ӫ S�p�`s���ƖL0%�lN�/Q������I�?�(j1�!�9T�9G�A��O�wHo^�٧1^w����f����{��G�%��є/�MN�Ÿ�u�]~I����F�P��]���̳ͤ:��O��&DK����o�@aAP��%",����K�j��|mÊ[
�DbD�r�����mh�4�E�bO��Ћ;���Iy�˻����pQԉ���́�=5~T
�u�I%E��=1�s(�bO%7�*h��ٚ�هi���|����##4��~�w��Vg2�%U���d{�P.�s�uL��F�8�k�L���U��^�I�%b� ��L������k���e���Hp)@
�kZ§�|�$i���O��5�4��X0=9�:��U�,�!��w��T����q�,�_�(�hpAv7D�cv�����|K4�y������f.>��]�7�-8-���3��.K ��h�Ǻp)�я��y�4RX;����ƓL�-W���%��m��^�J�B(,q>38a��e�!ٕV��zw^C'g�k���}&�zZ�ٰ~{�]~�
��I�n�[���ӊ��U�ȼ��le4���ci���C��)*1.tg�WA*{���Q&6��M6l�oӓ�}��>�(ܯ�$��c��˄�p��X�t��l��Q��b����]]Yյ�{���]/H��m}S\�e���c]�������N��i�{(�'`�P�+m���d.��E�jL���și�b�T�}�n�ij��Яvd���=���P���=*z��[�t9&�n������ǹ���	��9�J� �#�?X/`Bdt��b�z�Z]X�1�yѕ���'8l�))�ށ��O0W~Fo%��&�����D��7J��@�5^D7p��w�@E?�,��)i,K4�R�����!$J�V�xM�Ƣ� M��=���{ck��$�y�7odd�
�o�%�ν��Nu�
c�E��fz�İ���r�Ȱ(�u����|i�$�(|�/֧�!~.��#߂�����T�H�3�zSA�*�q���&��1�5�~��	 A-�`�/:`|�zb�L�d�9D��P�Oq����eЪ�/a�f(����aƝG��H���]]���Z�V�;"ЯEY��م�r� !�W�re��-����P��Q��Aھ�Vtݝމ�g ��rb�`�wtQ%h�NX��܇�))i��U������p�ʵ(�%�e��?g,"�����^�\�og���k0��Ϋ��uG�L�~4�f��Y��b�+��%X�)�V.�q_-�|A+�ol�8^��T����d�RXg!r�,�ݹ)z��
wx�F�d;-HE�vM=�i��*����B3AȜ-!Uc�J��ґ���v���#�����a�]���p�^�Yǚ�7;q�K�P��M��5�#m�Wa�֌r�C<�g�����]}�?p�(:E����L։�q�"�!NrW0˓��x.#:�,���ute���B�����r�T3�9	d�9�SF�1��p4�d��RU��J(��Mx���<��^��כd�Z߆�Z�n;#g�+��D���s��6�^SR�:���]dj[�#���F�G��r5Y�Ȯu��8�`.�i��4� �^&����
He[��W��aT��q`d�uD�=���g�j���F��6�g�E;�LE���%]h���r����%���&Q6���8��?���}嘲"��S��o#�[әw��"B;TT�VZwx���BX�ߢ�Gt�^4�N��wEQ(��ٽh50�2� ��
s64]�~@<?�L���4���|�%�B��lL��YG�\l_1�~�d�%�؅e��C�������C	
j���.�m��錼 k.�8�M���xf�V���IhЀ����{�Ez>.�]�a�~�:����F��8��O6Ϗ�z`�Z8������;WP7��t�.�]�j�[��hʗ�f3G����!�Q�6�|���C&�2�{���Y
ے����(�bH%�h�*�x'<��*��wΎ�C��ӻ[t\N�Z?��e�����A*����/ދ��bK������/
����.�t���~/����ʴ�1���,gR��ŋ�#�L�CFG~pڪ�a���0��s?���T�H$k";^ !�d�y}�:��OJ�����q>Z���R@M��=�x�Џ� s�SjŪ�[�١���&���2��st(q̫E�lmvt �y-��ל���t�meL�O��&���X��zM��Nv9lT�M�w8���"P��m�����U���x��XGQ����Y��F�!�����0��%��d9�~�č$,��0P{�%�c���>|�t����|�e�ӵA�/E��ߓ���/�`
酖�>Ne��g�Ɣ�^@�(֏�xS��O�ĭ�jH������5:����B���=nz�JV�oH�PFQ隔F�����ʱǌ��!P�`u[�.��?�,$�Br�ª,x��q�E�mzq@�W�n���7Gߝ���̘��}P*��A�ܴ@�d{F������(]�]���d�����૸�:�P�s�Wd$1Y㹳D�%Tt[����EXc�}j���_�wҨ~I٬�b�)}�QE©�w�-�<r�J�+���0.�oy��/R3���F���%mӍ*�b�2+�!:�%���tC�_�����ʠ�D׻Ni�K��f,9D�� o4]ى���g}2�S��ud~����?)�v��(�w�ŗ����9k�����%��S�cj�wJ��H�H���R�E��w��֞�8�A�t#����������պ�(3����pBk�`P�Z�3OV�A<�(�<EUÇO���f�R)"�BAg��%ئ�7/U�VÜ�������r�6\��D�a�/��M�df�ͽ���Ht�ǀχ�=�3��.c�~�a�3���#�X/�:7�S٥��NE���R@Z���*ȷ:ht�7p
�@��f;BL�� ���'+�ps=7{p��'�;��m��muK������Q��v�� t:a�Eu��T�@<���Ǚ�	�K�'�.7"~����t�e|��o�гbP>�bs#<�����G�;�����
�i`�ѩ���s�ܿ3��6}º�*U��4�l����g���_��71k�K�,uF�C����5�l�m7�Y;*F���p]��i`�����ڍ��!�d�ؖd8$k�ZO����hQ�^��1��I�YUm-^�t���C<��>���k��W�,ς��|�-[����N��K��I7ס��XS��`�Jְڕ���#�4��qDx�45���aǗ!lq��i�l���o�E׬��P<!jC���K�_���9�z�FtM�U����N(�J2b�N��x��L�FM�\A0D)����ST3�6߱��Eę�3�08�k��d����J)vd�=�ϰ̖��Z��W��π�7�СOſ�{)�|�_�~<�{�A/\��eJg�]���BD���=*�t�G�MY�"d�/<-��F��9�[V.B�ƅ�2�$�vc�v��>�-���x2{�_�Q
=i]�%�O[
����9����&-��눿�R���S�ث�$G
��"GA����xǜ��<��6*#BיL�u��ܧ$?���.��;�_>M��s6bH��ғR�Ń`.,�aӷ�+D~��R�[����6(����XX0\�D����٧�9v7�XMM�t;�^W�"��M��l�h�+�S���\h��Wb�����涭сn�P��hJ"� �9{C��ڣ�*-T�B0F-�t��Ō=^tL<��6�S���^j~�#���E�����d�o]�hs"ǒCDt�{)�����!�rcK�^]�Y}���H��WS�*Bc�o�pҷ��p���6�ջ�q���d.���&Ң{�!��<��&���y��
����U�C��O�CM��UAxoSֈ���6�+E�nW��?���d�'�fh����j+����I5tV��&{w!�y+���bXY�HS�J_o ��T��Zz�����J=BXH�F
�X��5�(�j�h���~�5w>lZ������,���t�F(8�� ���g�,�ؤ�EkI�yqm�h���Ld���hv���FC�H��N���d��DA��`Q�~����I������\�I��
��������!�=�2��)���/aj(��}��me�1�
w{GH��^�aD�5־r�M��
�_rp<_�a|�\�_�}�儊�������৸#�6��E!1dM��im�s0���2mt�����꓂��?�,0Erh�5�F*��W-4j��j�A=�,!y�����IJ��i�t� ���f�p�?~Q�5�0AU���h�DΠ�m��,��m�o�*i��h"�sx��ln.�k��l<w$��t�i0�	��U2�8�l�mj����dی�iz���V�\���Zqq�LK�/Y��]j���!=:��� .�c�u��:^<�� ���r���f������4�2p��l�H�oZZLĦ��l���SAD{ 4dʯ<>.�DA���Med�̓7rW��R&��Xz1�7�ƀ9���j�}!�Ή�l$���̬�\kWV'���ܢ:zD�邭'^^��_�8��"줙	��N�`a�Cm�'0Nn�?i��%�!=�ޣ#:9���A�Nv�0��=d;�1+�[��u��l7͕Ϙ��g1%�U^���M����a]UԽ�2j���W�8@^�yb���QX^�/���V�[���|���p��l,wm� �u��A�)?ˤ�r���l�l����]͛"Y�Q ����a��y�W&y�$�g�[��1q>cJ�/z���ے._�|ǐ��P��%����m*��h져{@t����uH��z]�q�2NJT�~��tiQ�s�5=�M7#�y�(��*|�Fk����}�O�[6{'$� �(�Mq�X?��ǝa�����3�i��[��/�zF��������%5�c��%�Ơ�_��==�7]���X���o��m�zҒ�	E�&Z�Z�& �h�v����mp=#�^d'&���Gѽ ǬQz�Z��Պ�Ss�W���vKĭ���u�4�2��Lz�d���,���簮A4K:f-��n�Y��	��z�C|�j9@�Ֆ{G�A�ǫ�fq���,5Hi6�;�PX�Z=��q�C�uqe=��t���h��:�z�����6�����A"�~Owh�r3����{����Dgw�ϣIF�K��E=���2�wW�4��D�M^
�68���x��>)�[�d��R�M��'�����n��`��⏘L}������|tm77[!�ݒ��BsU�7��L���0�%ν���w�Q8��ԏO�k�C��_���%>�
Ұw��Aup[UA�H��k���Ñ���&6Ͷ���̮��.P.�¹��&ܫ�S���9�ZtI[�+�S�ߥ6�V:E���o��z8�&}&���sP����}�6��!�"^��"���p�X��v%�D\�>�J�t�!�>�9��桶��K�Ŝ{�^~�D��J�-W�f�*4�//�_�Rl@���@��~B4:�;lR�-f B�e`N�o�宇44,��S�/`Ĩh?![�5�[)3
BN�m"y��&�L4�+0�m�7[�P;�˅��<���@!�~<����_��#;-QN�:��X��.s����	�ȧ^��0&Y�_^0BF1+��%�-�w+�r�l+.,�?x!��X��-�'�n 9hKo1�x��v?X��MM����׳��o�Z\o�ᒸ~�S��$0�a�`2_#�ܘ�.�;Ǹx��ø#�9v��Ms ��(v:5�PܾM��ntI9�i�C��� �Ԣ�'��-R��b�p9����s��/���ALoF�	B��u-�*�jG���%OS�ۊ�S��ԛ���i�w����b��_��CF�8��OԘ��E���K��匙"�<���%ŗ\��@��_L��"'�h(e#_yI�VOKZ� +3%���ɻ�B�v'��'�m��H+����%=>�z���X�D�)f$�8�*[��oȝ���MoAks~$,Dt��W�x�d����%b0�5w���?SXP;z�7�͟�ٸ��H��~��"$n{���G��|J���̄CÂa�=C���Aɗ	�����8�ެ��5��.�.~��ܱne�n��(��a����bf<vL�Z��Ьn�HS`c�N'�8ŔfH5�67Y�BP���h�� 6�+V3}���l� 6�u�j�e��&�UڣE�:`3��zX��*��
1R�����:�G$eU�P�y�~��R�v�(��C�J��f@�B��MW�=��lL�B���g�{zQ䩃�ZV9]!��Ө2;֧��A;���nXJ*�̓�p7*�-�lO��m]I� Z%)1�vǓ�_@eWP��&���G���E�b�,)���
���O�������0��++��!��+�@Ȅ�s�]���.���!$�%^���}���Ve`yG��l̩=�o��ǎ��"�|N2�,�������q�� �bb$]�%�1ҕu�� ��7R�yK����<fP��?���~�!Rv����|$+�y�:V�kH�!�rWj�-Ό��YL��]~`��gKTmU;@�J�h�ӳ�I(]*L�0sp\h����81����麜$<�V��M�����$����gC����`ˡ(�$��N�?�b�0���z���
�"D?��>W�#�Ǩk�6� �N��h��%�X>�u��'�R�F�-B��=�����2�	@��ĭXל�j��̜�Z=IJ�e�R�	�pl5{�	��1�e3V��H���'�r�w8����v鯴�Ή�_,74+D��#�Yq��`Q����*wNFCN�Z�b�� ҜS�Ê�*I%�N��g:��	&+��'������Г��!zi�e�T3�m�$+.��^p�����I���+?!�|3�����X�z���4t7����/�i��[%��q�!�3�z=�_�G}��~\�pZ�4�lrb�s�.�f|C'����Î���N`
Ѝj-� �V)��$K ۞�����FF�a����	d��@)8�!W�u>öy�K �/qV찜�
�C�1-qn#fmΛNp
��KBr�������:�iDA�/Y��:�3�(O����ɱ�n ��)�cE���Cf�3v�d�R�+��6��y��v�)���)e ؍�2�$�z`E!�v(n� ��:Kt�ѭ/T^�e۳ت	9Ri��y�;�<��C+!�[~C�82nBj�[��c��E�B�jFk���;-PZ��PgA��L#8@�x�! �̊�8�_��nǻ�6�_�|Z�l�#��T
iq��3t�*I+( S�~u�|�B�v�f�	L�)���J�{��ﴧ:�,�iapZ�j�S��X�4�B8�;LH5��k�ĤeL�~��ƖMڳfs�'���%���6v�._��\sKʀm����iex�>!S�$�W�On�֡�ܔ-2|~��P��	 D��dq�S!,��l/t�Z��]t�Wa��*�|����^�f��T�p)����t�Ue�TP�ܕ��2�VNdr�PL����r$����������������h���0��XcAei쐛&^���v�B�G�$��@�$�$�������m�<��cœ�y�i\�)�5#�<"��%q��0�z�[��}���6PB8\;OX�qR� 7V&�A��s�?������HP@/�(��7q�=�q�oiW�'_^�b�~JsL�YV���o���Ā`|�iQ����@ǈҘ�]�	�)(���c���7~�h�d�b�sI!�6�M�Ka��N��-��d��*�	�F<�g��p/�$9����r�nЙ�I�^��Ť��//�����0=����������4@z<<�@Z������a�� �}�V[���吔�W�0��'Z���|��j0��d����<���� �����-Z=VR؝��w� ǭ�y�V�CU�',ȃ�p���s�5�h�-5��R�
�$�b��e��%�X��Q��7e�M*N./��&��l�4<��J����mxĈ�L����.r��ހ�Uf�����N)�[�%z�6�B;�y����;�R+��!c�ۜ}s�|�8}Ȳ%b'�Ҙ���Ϻ�-
��˴a��Q+��xO&���I�%x?��'����X吽(�$�� 017����XqZ�#V���b!�Q��M�5�p��vv&��$�n���E�<l�C�B1E�0Y4� �����,S����J�Yw��6^{9�]���p.fSW!�U��0�y�E�ױ�,ix(����,�c+����9|m��`O#����<p	^����<q��8�@~�|.��M<�ݽ���l��Lq���@6�-l���{^��u�k�%}ǀ_�j�-U�=Q^&�Ƕ�ޟR�R��`^n�w�G`8�F�b���;���M.�e\���]XkCjC��XB�wM�?f��RYjZzVk51�(�x>��2S���W���'���i�Ȯu�I�@AkE(m�|,��jU�Qyޖ'��"�I׊��8W�\GUY�6��Q�D�
4K����|g��8�-����6D��d������"�6�1�եB��Υ��z�@ҏ_1�B�'����<zT��j^&��k�X+$dm�/H��%��&���M�ؔ'��J�"��G����K�������0ӻ��[��d^�����Z4H��Ը�7�ӿ$��L
�󗑏�+��
�����竞�v�w�ڬ=�z�~~��}�O��F�m��+�EA�g&N�K���1��K>���\͙��[C�c�Y��g�Y��2�}�@�RBo��اG�zS��Q��	Eܐ�#ߎe�f��1��7�%��'�������C�m;S(��P� LJ��&2P��.�uy�r���	jb�%"�Z߅�3��l�;��;�h�������#ѓ�c�b��t}�4	ғs�	M"�ZX��
��V��_��͎���Gm�C�f�V$i�Rq��Н̥��X�q�당��M@%_hiȢy�F�z �(<oA�V�����0��E%��`ڳ��<	*�N���Y�y@w_��1��7���(r�N=���q<�\T #l���'�L_s'B�2���}WL������ǀЙ�R0��)ܯM�^�����b�k�a2-��"
J���&_ �V d8x��!���˟�,�9�g��#-�ݟ��b�F����M��u����_J���c��v������6��o� �?��2inȐx^4��_i�X@�L��:8�)�2��k�r���q[G�P~J s� �}khz�����l+��%{DV�N�f���l�m�c��>��������r5E �}����G2g�������k3������&0�n]hH�ުH���ʰ��דeC��-���/��b�ҙ�[p�Z:�q?
�{y�c�]��	u����~�KC؍�!X�HB����e�����/��-p<�.��1���`�ƣuR�t�1�"���}(�ik����fZW��qV?��[�k�+QM]���=-���m��&X�[���AeT[{���@7?���^)#��Ǐ�$�ͫU<�ຈ��P��U8�m;�a�WxJ��;j�![���$V^���Nu��ьdkw�(Cۥf�m���ӀN���@�ٵ��`�t`~1���L}U_5�]:1��[%~� �Ҹ��F�(�<�����Ƌʋ��)��N�����|Zĸ.���LGP��ο�>��A�V�+�|�m;o~�s�<�I��wu�F�a������:�$COTtE'��|�X�Z�Lꑧ���P)���J�/B����}�-��Y����|��ڔW0�w[���� #��}�&^BǍR��J�J:�3�C@��)�-���b��Kq[��ǵ�Jx��Vd�;�F��>��Nqn�[��0�P�?Ǚ0��,�����5�,W#{����(��B�mv
��ﶂgh�B��K>�\�9���Z_k��a/K�po�Ep�����`:��8R�a��E��]�h��;��m���_�'��	��+xէj���^4�B4M3ç_<m���t���R!��	��_$�	w h��_2Ļ�ѭ�mːNj�g8"���}��m
�J莋�9q�#jA�v���UY��3��wah3[1���ԋ�B���<VT-Xs|x����\;����{A�7�CY�}�@0�V�"=����k���qXvf����mjtV>�'s'@�覦���n�y��-ɒ��<v��u|�Հ��Ac 8�dП1��h|˛PC"���M���$x�]�7��E��'*NŲ�!d�wV~U�����J��.���{l؅�yE�%4�	N�=;���F S����|O/6��`Oo�@�(~)PWR��L�v�"��O�@#�W��=j^�ZTw��	dn�����N1���b�kR��b����	���1O�u���Q�Ŝq�3�Nt5[��P��l޴�[�أ���(BҔ���o�2=�7 �Ȃ�V�OP�o�Oڴ������g�]����Ω��B��T_ �T�zB=�Ý�UrfD~}���V�4f�S���8�D� ��v+���k��
�ЅAH*,+~46���k���������E����Q]+<̉'�=�� �t�,��������w��;�-�	Q:&u���\��#��O֑��@�}';���>M�smQCۜ6i��:\o-雗	���zV��-\v���|����o���1����^[6Q�փӻ����#��ρ�9���ڝ�K����x���A\�V#�k���P�ʪ+�"�

��:�a��Q��2�Q69V~VA�� 1F�"?$�w��
�i ۸I�`�)���y�ww�A��t�����~�S��l��n5e��5 �t�X�����{�m�����M�a��>t,�P>ܢ��X��-v����������N�f���dj����lh���a!/O�V)�uӈ�?���v���B.���mɫf��ē4�=Z�H�-{���a	ӵ�m���9��JX���-4lմ�4��g���S�zA��X^��0��׽Y3�:��1��+���ݳ{�� ����G��5ɽ�ՙ<}\��t���O��E��1{��,����F�¿`H�c{�A��F$+y�0��KI��ۀ��v�|� �Ǚ���r�_�:<�"$C;�6�¬�E&8dz(]Nz7:v�[�椅�?�
TU�Hb�"j�-��Uih��|Kc�o}nzG�ņ��,7���>���ꉼ��=��@囲( ��id��?��y��n�V��N�LC���O瞖 ��O�M.5-Y:�9O�]	�Co'f2�P>��E���Z�?���	2 ��D
�EX��������'�T ��(�圍@���HBu��m	� ���\%������3����"�2�\��ؿ�G�hL��*9Qp�0��u�!%��Lf4����\�h1�s�>���5c@�a-�$�0*w�$�p4��`�KR�����:���n�ո�����3���j1�ȏw� z�����I�k)�;��Q���f��u��tRo�G���|�?���)gpp����0�F��m�'h���[ytce�V+"y� ��������m���!�旭}�w��ܑxW�@�-G�oh{�� ��T���g${�_��&�qZ����մ��=�-���K& �
{��Qq�~��?^�G#�FĠq�����=�!�/�C-y�S|vռ�$�ۆ�Ve ���OuZ���|R}Ȑ�9��z?�n]�iJ��}M���'Lu])��&��hr[�x���-�o�!ey����D�8�&J�w*u�$�8��`<�K9�I�;�_j9�tB
�L?2����5�.��4���3ka~	VZ#�fe�Ӿ����k`\ܕ�`�\�QH��YP���f��DWiT���`M�P��!%p�,���ÜW �q-�~��v	��h�vav�Y��A��ڻ����DQ4��tq���-�a�khZ+	~r�գ������>;^9�Q���1�T1�
#��/ȟ�������ɏ`�J���hܜm�?�aa"5�`���V��Ѩ�W`9�P%�m�*�mu9!S;�6�h�#�WК^_���<�[[��,����|8\���r�}��i<je���%χA��<�@z�7c��/��.�po�E-`�|K��2��inZ[�����o"�V���=���}�z>Ih�	t�^]��x��#X��+mt(-�ޞ^�#B��U�*%5S�g���V�4j�Q66���*Sj��,Ȍb�l�$[Mp_�$�������F�쫲���Z�Ö���&��� 6D�G2�$E�0��r~4C��c/�`�^����Z�4����l��;a�M��ۃ���V"e�j!���`<�)�IW�*��2��ql��x��D����CU3�*_��v.�_ܹ�!X����_��[SH \v)5ң����n>Շ<��Z�;l4*NR��y�m
Q����#ɘ=�v�4P��i�f� ��N3�C6���l�u7�E��;x�i%2����*W&� �cz��S\W�0%��!��5�K��/�*]Vo�:͡b��Ӭ2��ʱ)L��d��>�F��IwN�1w���aת�MT�i��yӶ0����v�	�t�Y�4����Pw�LN�l�i��`�h��=��� ���(�_��l(٘����k��$�;�s�E�V�����ɪX�\9�����9�u����@��AM<�l�H" 2춆��Yfp��
�����xl��Y�Av�;�%7�]ʧѶM�{r,?dDt�3x���漑4����!mq�_�$������n�:�Z5�����SAMT�@���f�|x"�E�}��Cerz1���V3��gN�4.�E�7,/��
�y��	�L��
c�~q8��B�Ay>*O���V `@M�Ś\!��v����[�R�T�Q����Fg������)��l:k5�*�vUX��MaK� �3tA�Ȍq��uĪ���Lo�l`0�l{R���4YO��6d���DU{T�9�h	��L��OJ�o҄:oӛ��U4"eI�B� �1Q�؂GWm	�;����M� S�����`��,��g:G� �Y��C'��v��G J�N{�o��wv	,Hm��$��e,��e.0V=��������0A8��H`�����ZS�3뭕��!��� �K���<�q\�I�Wl͝��te��c��]q�?)bY���f޽i�[nQ���� T}�jD���ϊ��I�=���8�odF���/N�P�=�-<O�dM��Q�+�n�.2	?�f�D��Yݣ��6�@/��8b���d[E�����.d�_���Hm�P���:�jl�TɒM4�;:�B[�ʚ�7�2����pH��e'$!Z�y���D�5?�塬�!����4cU7
5<T�)��v��Q���>������'���ٳ��UO������Q	@�ذ�N��f�	(�qk?��Щ�������2�1k"��%�ƣ��>%|QFj:�/_�N�\=$��:�A�B�7�B4G1!nP&r����g�B�[�W�
�$�C ��Y�����2�݋XN��w���p�K�M�#�����������DI�W����Hj��H۽ߋ�5�GL� fѰ�U���g��i���B}�5�Ӛ�%N"1�����M��:5���޻0�ȏ�A�� �An`�0t��u#��