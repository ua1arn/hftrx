��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω����	8�;'N[��I�]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPy�����h���!�}�1�:�Ω����	8�;'N[��I�]P*m����)O��Ξ4�"�\�� ���K�O�{��׮���^�ן��A�ߙc\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��"O��Ą��J��]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�Kwz��
����J��$mm4rz��x�@@m	G��{cB�38���E���2O��'HY-٥��2*�D���J7"2�i�$�;Z ���������	x]̍��;��7�I��"8YdK�o����Oh5��&}Xa��gR�ca������pN�Wu��w)�S��X3����~篟|��ᕧSt ��[֊��Jџ�_�v%䆘[m�~R���\D�	m�!=�y����h�}�)���32�)���K��OC���N^o?�M��;]���i͹�9 ���t��%���&Oǀ�Һ�3{����V���	x]�<���eQ���X��\���|�@c���Կ�:�%n��e�ι̕��R)U�~�O���`Y�5���=�zX4P?�o��ľ��UW��͌Tfu��w)�S �J���vy7��Mv�9�h�s����b�z�Y8�:r&@�	��Ϸ)�����V\~{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�T�`�7?�\��4�/�I����D;�~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/�R����+��T��D[I'�p\���nEA�ܵ�j8�y�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcJe`xҖ3Ӫ�1?)�Cu��şo��q����R�_8�%���7���%%�xg��ۺ�D�U���&��,� A���W�F�ݸ��]ds�lOLH����DK�$s��?xA4��?�d���&�p�m~|�֟j��?q��N���%�5<{��T�O���6���\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�V�
]sNJ�}�+�r1D��y;�L���9�D_�3���U_�+X�p^'�&��5F:	��Q$n�tiW<���ubr�N���,��o���&W�Gj�x��^�%�|�oT�C@��AO}$|~�K��������� 2�D쉽�3CN>�4�
��}�`wKݷ�F">[P�9�g���Iv�䃨c^��Q/)�EY[��g6�w��U�N�>@�%� �,+��T��D[I'�p\���nEA�Dx 1�"(8<�V�Zs˿�}w��^z[��K�j��c�s��v?�%�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��W����&Q�Vdĳ���;t>
r?����x�fc��7z=���x������<��.�`�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�ؿ2�%��ĕT�u |��Gj�x�륗YgYM�w$���K���6O���d�Uf�揆0�бԧ2N��n���?���^�,ԯ���gnņ��#�b��~�26��\_XUfm>��x�ZWEב.`�Z�����èV$ Hl�]���'�PD��q{�).+�b��!qq�i7N�_��@��s���՝�6Ǻg��������:=H��Alϊ�$uEN4������&G�/��@���{j��ț��?	�MG`�g���j"<�i(��M��g%MG`�g��Q,����	~vT���f|O`�� \)޼QE1�D�Y7#iO��(O�T�}Dq�f��5ߧE4��HN��R���מu��� �H�0��
�y�"�V��5M��z�o�OP����z,7�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��h�>d�q/@�� "�s��?y]���4.\�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開<u��R��0�z}�J�T_��2��ۦ� ~�p�ޒ֙f���d�X�VM�����a�"y�ӓ���&D�H��hC$?���;���EWr��&�}'7�ܥ��2�o�{e����ś���k� ��b�FP&� ��Bo	��%��r��Y��d庒��� л��l�R�"h����m� v����5E�ۼA�}��ֱ�q�����)���p౳�#�^:��L��XmΘ�# ��b�FP&���x�Źx��4�o�rޡ����u>��uL-���%K��ͪM$յ[+8�V>�V����,��b�z'hۉ)�禫����#^���,�x�<��V5+��:�M{�����q��L/L������([ˊ�����|#HK��&첝挅0����A�.1tSjv�֭�h��Ou��WP���� #i�_�/i����&�}'T��0aȜ�}Dq�f��#^���,�x�<���ݚ�Н�[J@&�4����/M������_r��ݚ�Н�V>�V����,��b�z'hۉ)�禫����	��x��ݚ�Н�V>�V���^�w"Cj����*��Q�ܬ�:�B�'��a�q�M'�y�?W�k �b�[�gMh�fĉ>99��A0ok�?�JY�)�Y`��jD4�B�h,d��Z�!�f^ �W>���ĕT�u |�T���u�ܙq}ĕ�!��(�
@��^���3�}@��9�ڮW��J�	^�M����A��}�9S���;xI|$���"�|�E+��T��D[I'�p\���nEAv6�	l�