��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�LZ*IV���^������0K_[��e�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k��O��ڴ���WЋ��I�?g�f�ja1�n�[�c�/�O��?�;��XC�V���E<v��b1Ø^���#K���lӧIA�a�V��R��tv�Τ���i�wJ�'�دv)h�V~�$v�p��"}�v\-8�������>�`)���a��rl�ʩ{�Bf��� ��|4�VDG+�������X".��>��'��E����F�Rm�I�|^�Q�;(1Z �bRw�����IL�+�{Dr[��	�� '�T�������3�f�_��ic��H9�~r�_���TF_���TF_���TF�ձ��y_���TF�ձ��y�h4�h��*����~�{4�a�
��!�`�(i34�a�
��!�`�(i34�a�
��!�`�(i3��g��~�G���s��4A��a_8|4A��a_8|��K{l�+~��c�'��K{l�+ ���M���f�}.#3����Fz�!�`�(i3E�V�.\*�!�`�(i3!�`�(i3!�`�(i3h��ٌ��!�`�(i3�+���4���Fz�!�`�(i3!�`�(i3ef�m�5����Fz�!�`�(i3!�`�(i3!�`�(i3,��L���!�`�(i3!�`�(i3!�`�(i3Kp(����Q#�y�&(���B��|�(����5���I�zI.��1��b־���1N<��;���u��w)�S��X3����~篟|��
O�:��t����;r8�:r&@1�+Q�<��d���L!ۤՀ/Q9*سBK-����s~�j1���u��w)�S��X3�����@��."�;r|@�b�؃��em�J�Й�m��JNu���]�ߏ��P�umSe��S�2�:,�nr#�9l$�/P��pO�c�c�ENk�lAc>b�G��8̀@��k.�"SӠ�|&��c���m�Rܙ#l�%q�M�4�}�����r�N�Þ��t�U�PD@��k.͇�@�L�v���0�Rc=���T�1�\�^6uk��~1f��t�jPP�
� �AH����e��'�Wا[~�l]ǜ�����] ��F@�4%���D�Pfc����2P����/�"��< ���X�M+��tc��P9P��`�.�D���J7"Xv�oʬ��
r:�����u��w)�S-!�����c�J�M=�r�����|m�nyZȕ8�:r&@f����:dD;CBs(IkT˱ �Y�p�3c!��h@��u���
|H?���v��E�?�Y��}7]4Qbt�_�݆��5R���[�ޛ��g����R�u��w)�Sl���-�edc�J�M=�2��&�	��1�`�a8�:r&@�G	���su�]bu̎x4�J��|���>�
� �AH���CdZ�G�u� �(�a�b<UӨ�����"v��J�Й�m�a�|goS3������~��Y��6����uS �����t0+zW��D-i���w��#��D�?F��,7�j�2>����.z⥩'kr��{ib�c���I����uS ����ߩ��,j� c��(�U����	x]��Y'��G]c�J�M=
��%j�D���-)8�:r&@9����DY�Ԕ/h2�Ժa6��(�����~��0��-�y�xUq�}���hv�(��z�j�#H�Z�T�+?3�l����ە� � ��|��e1����� a�;qPƵp��
� �AH�W���,2w���$�cUY��p�5NJ��f���F@�4%��]��N�"�<�/���;c n�b
� �AH� K�`A���vJ�^ <.���f�'�X�׼J�Й�m��C��ߊk'�4+.���`uI�[l٧cJ�^j�u��w)�S�5� �7��Mv�9*���f��^(��f�)y�8�:r&@��=��$얃�rb2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEA�����G��KJ(𬍝��;{g�P�r�|A�־���1��}�����b���q���1�:�Ω�S�T�;Ϗk[�^��_�6A�7Oq�@5�.ߖ�g��o�4��?��d��q�G�+��T��/o��إ�8p	�rh5���Z=%��dÂ��t�iZ]XF�������̘�иܖ��Q�P���O ���3�ҺIÙ=�H*.�PS�������Dɵ�p�AJ�e�$�� nU�IÙ=�HF���m¡p~z�r,����� ���3�ҺIÙ=�H*.�PS���ct�:��RE��]n�� ���3�ҺIÙ=�H<z,Ҽ&�כ��p܏�<
DN��Q�^�y�zL͊�q���Vǃ����B�6�N@���k���E����F�'n�^0o4M,�����t������ݪ�򈟆�������\�vņ	N�1�.�]V�H7'�5�}�]���!�`�(i3x�]�V���	�?�ki%�7%1�e)s 3�:��)�[���6"�,�>E��4];ˍH�,t����t�i�lK�I<��fҾ��9��ЂDa��(o��0��7Y%T��BPe.��xu	�>��l%i�-�M�g����!�`�(i3v�ј�"��Z鎬����F�71�B��>c��?�"�,�>E����-��%Mό���.�q�\E��0�����?x��#��]����������ݹ�0�����иܖ��+V.���w¹��<d���lC��U�T�\ �͹g}|�H� 7�J�[&e�l�����-��%Mm�jp=�>��o�
�v�ξ������eiy|��!k�R�^Ƒ����"X��[��Q[R�72W���R0L�>��0�]2�y�Z鎬����
C��8q��f�kN�ı���}J�|���|���O�.��_$��Y�7#�xI��W��_�ړ8���/�I<��f��tN2s���(����5���I�zI.��1��b־���1������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©��'w��
�f��]�/V��Xc�u:�^Y(��]�/(f�|��*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P�|h{�T��`�)�	�%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��Vx�%L��W��_�ړ8���/����RY��0!S�,��ш�A3�(N��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���_U)�<�&#R�^Ƒ����"X��[��Q[R�7����n9읣_--���g�vh�1�WpH7���
I@1�ؠ&���Z02��`�z��GZ>.�0�i�ܰAb!��u�mj�B��Vhs5e�U�Ͱ��Le�2l��4��a��se�ξ������ei4����/����DP֞ �����KE ���1P�]�׼�a�r��AR1<]Q�I����q��� U����z~�����~�
_g��c����o����W0i��^&$��}�����]�w�r��VYW\y]/�qFtԸ�7����|�����-���V�T_��p��כ��pܚ����U�Op�m~|��4��ݬ��0M�/�s����Op�ե[?M-��6(uU����z~-� �lZ����$�1�=z�>���@�<[n^/��u�h踫g(�r� k�|6�8����^��L�de��y]/�qF��6��	���`y���h}Nw���U�m#j[3���w�@V�/�˟��7<���������	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8��L���N@�/�M�9���{p7�j�pܔp�l
d�R�.��On��M��ҹf�f3'i3�|)sՀ�/V����!�`�(i3���^��=z�>����ep�G;w���w��l��ML�f���|����OxtX+�Y�G��"j:}��M�+����ei�}�"Io?�?��A�^kAO��t�+���LQ���"X��[��Q[R�7��iM��*����6*�Gc_����+�˂߮<u�4�!>I�W��^�����f��|�F7�_��O����2ا@����\+>���y߼
�d�5�a��3�#ң��}�o��>n��rs�i�a�}Q��C�q��2!K���ž�N��� <&�M#'���Xwd�n]N�hC$?���;���EWr����Ly��Y�{'%s��v�9˞�P�)��j��`y�����n4s1�h�9�*�?�j+c�<�ܿm.��ٯ�<�e��BF�R�\<۳��Z�^��� K�bXox��'ѧ�#O&GV�z�<���Ŝ�0�Du�d��/���
.`��}φ��R%m�Rs��R���:K=c�CuV��B��K��3&%��^[���F��O�ЂDa��(W)5S�7KnZm`�x����Cҷ��e��߬}u1u?�:�H�ܷ1ŭM�,E4SG���Z����� h�ҩ��i7N�_��
H�(1���P]	G&N���k;Q?M8�f2o|���P��3 �n�R�]c�����u^��󀋄�g���W0�]��e|)0� ��(nW�'{w#/ B7�%M��4f�x #^�9n��,�J��/3o�U�r*A&-�Ri֭�h��O�\@Ui�-ƍ2���lķu��A�0�Ή*��a��71�FHN��R��bP�63Z�t��\�Ж ���-3��q�l;1�U������Eo"'N�q�ȓ�iӚ/Syb3kP8{���@��u��_�����d�J��:����(Y��:���R'cf���³5��&l�����#W�U��ظ�d���!i�/��@��C�G����]'\gWg��	�Z�kfc��2���8[�����(����<m�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�?V��j�c>ݣK�6<o�k��G<Y�dN�<@Iv��nt=:��:5A��p�B�'��a� 7�J�[|�m�ߕ�E�g�������(ӈ���m�r����!�`�(i3�k��M��߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv��!�`�(i3y�}�6f&rG��Hb� h�ҩ�!�`�(i3?KYC'v���ʗ�%���S�*(�����Ə!�w(�y?!�`�(i3��nސ��3���w�@V�  ����'mj�B��V3�����n!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��φ��<�6���%5)RHN��R��?�d���&����yϔUw�R���y���,!��%.gW>�a�ut�0o��F�5(��~�q��a+��bc�n7�}�!��?KYC'v���NE!/ ,��rQ�i=�d�ЈH����@�/�M�=t�z 7�J�[4���0���V��	��y&Qe�}�!_aP6r��$����i7N�_�Ar��� ��иܖ��A�.u�r;��|B?,
�H {��u��]'\gWg��	�Z�kfc��2���8���8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�7�A��\RE�g�������(ӈ���m�r����̢k���"��w6�0��ɗ��zi#Y)M���Fe���2+m�7m�T��Ʈ+ˀa��z��2�,�s�Yls��8��GM2�]�<�!�`�(i3��#
<�(z.Ю;�Ƴ0��atN�s��S�+��ׇӭ��V�Ո��Ú�'nB��!���c�A�L'0#P�O�Rfł��kS�*;q��
�7Cv��L�*dgN;�r��H�?X���V4&v��؄aX�
�:qEp�q�?^�V!�`�(i3��4-劽51�X�c�rs�i� S�xSVe�W�6?���_--���g|�m�ߕ���s���OgE�s@�@�/�M�[=՗Rz5�(��&�����%>�rGO�D mWN!�`�(i3=��,���H9a�Fc��Rfł��kS�*;q��
�7Cv��L�*dgN;�r��H�?X���V4&��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M0���w�����,�ǰ���!�Ab�����n�-�IZ��R'cf��w���Q��O�بeD�Iћ���ڀS��d���!i���+�^��BY�B<C�.���pD9|�
�wFlE� ��*�n�'���"/blU�5��Dz��6|4E98�5�O�%E#P`6���ҹ"��s��?%ww��Q��ǺΕ�=Y��~K?�d���&��ݚ�Н���hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�����o�aq����1S�Д_9[�l��a+Ĳ
�),��Tt�j� �"�m���rwӷ9J�E[�l��a+Ĳ
�),�5C��-��"�m���r!|�α+I��)���W�w��fD��TA��w���j�8Oqҹ"��s�wP�>Q��ǺΕod'ٙ� �z�:Y���J��:����SƏw0��C�ݥc&���XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���Zt%��m&<�P8��PS~B;�T��Q׭n�L���/=9��9����C.�L:,��i���A��;b�-�2�V��	��y�9z�Q��S��}Dq�f�Hg�'/�F(+� �e���5*s6=��GZ>.�0'j�j�Jy?�d���&��ݚ�Н���hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�����o�aq����1>� {�}���my$�N��o�/���;fĉ>99��;��|B3���Hρ��~�_�=%䟳��L� *NK��阬иܖ����S�f>x�:	�W+��W�FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���r!|�α+SƏw0��C�ݥc&�̢����{_8�Y��=�}�Vݨ��}Dq�f�����,�ǰO8l5��E�i�m}66j�"Hs0vZ��ҹ0�(j��0�S��q�;��3O/tկ�oȺf��Ҧ��>!s?�d���&��@��v{�G2�e��b�uX�R୊MEφ��<�6�@a� ��fFMqlgC>��Ӛ��S�J\7~�8�r\���1 ��ޣM��;�jmT�#bs��2[�a��o���H�RtV�^FkH��۟�z��n�*�&�v��K7͍��|��W&":�ݚ�Н�!q��V���<	s/����AIe��0�U+�qbp@�!�`�(i3����g�Z��3��a���!@�f")u��r��;�jmT�#�,l����M?��y�!�`�(i3�Zj���
�%q�>��8�>r&���c
� �ƚ�-����!�`�(i3FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+!�`�(i3!q��V���<	s/.�Ss�g��+˘\5���jmY�VS���g�n�{�6�e
��>�i�g��+˘\5���jmY��X"e_�4�{�6�em�;���!�`�(i3�k��^�1.aIC:L{0w����u���ei�@�ܫ՞�� h�ҩ�!�`�(i3��hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�!�`�(i3U�~�vmȋ��OY'���c���鿋�E~��k}����/]P�����+���LQ��:5A��p
�:qEpA� ��_��5X���иܖ����Sp��;�{��!�`�(i3Zt%��m&<�P8��PS~�Dn��i�Q׭n�L���/=9j���)��Q��\@
��:�)�<�����⪂!t-�u	D�&���A3�Q��\@
����G3҇
!�`�(i3SƏw0��C�ݥc&�̢����{_8�Y��=�}�Vݨ��}Dq�f�՝� s�#���k$ !�`�(i3��hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]��}Dq�f�!�`�(i3U�~�vmȋ��OY'�E�g�������(ӈ���m�r����!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹�%G��^���j�VD"q��_N��.�g3Z-:S�4��Y�Y8��t���'!2t썿����`�φ��<�6�@a� ���N���������y��o��7�;�jmT�#bs��2[�a��o���H�RtV�^����o�aZⓞ��mdN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'����u��r��Zt%��m&<��3�H[ރ��Ŋ5�m��P8��PS~��\���
�C�ݥc&���2�!�,�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�� �ѕC?"_U�In��u����,�ǰ�QCT�"����Vx`���5�� gWVbT+踫g(�r�2�������l혡˩��H�V�����,u�x{��̷_��yC��S8����ڝ�̗g�Nri ��/z*x�n;��|B�%5[��xx�FX���v�\�b�U4��\w��˪?�-���ei�^�̷ؠJ��:����}V�)c�`j�Txk^��]��3R��������Vo[���˚����Z���2��}�������Ə�m1�ؓ� ,��rQ3���w�@VeX�P�+$r�t�}iV��	��y�� �P�qN#?
]w<�h��R��e�j�Txk^�a���~6�z�����ϲ��Vo[���˚����Z�ם�.J7h��r��H�v@W��}�������D3���w�@V��B|_��j$r�t�}iV��	��y�� �P�qNy�WE~�YV��	��y�2B��$X|,�E_�CR��L(q_҂T�q�w���Q��O�بeD�Iћ���ڀS��d���!i��x��=;Y�ۺ�Ub�!�V��u��i�_:���5�%]����8�B���ow_;O
�J��:����{k�h�+*J�X�$��+�nj�a�0r�uzZa�U2X��������,�ǰ�������� 7�G�Yw�R���yWp�K#J���.�U �3Ah	)ޟ�I.��^�