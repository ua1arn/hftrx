��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p ��%Dr��hu9���c*�?�m��������$h���Pjn�N�P6ĳ��@�o����`~�ۙڰ\2�a��-��jfPG�����B,t���Y�!��/a'���<��?�SvWIo��u���Jg�����uE��K��"�V<��R���h|��Eя6n��؉%�����Ez���\�L�^ߪi}�>�;��:5��#���=R��f%��ѯ���+^�i�M��kO�����AX��hة��Ԍ+)��N�W5g��i�H8��=�T@������)�s�]�nT��4sU��'
wRs�1�ʪ2�<�{0-���K���M�0��Ƅ�H@�� �]t����cHԪ;��w%ڛ�p�D��X�;����-8�93EM�c���G��T@�� ��},�V��N���	�_���� ج�pT `KJ���L{�t+���ԄK���
��_� ��C1O�@�B���
%��"?�Gm����d?�:g�%�ѱ����vM
/�İ'qRd���.�I�n�����dk���06B'=���u�v�<������w�,2��niG�M����>�&�|�A�e2�w��D����&ib����oY��
й��,�����YJ��#c
4���T��"�z��6å7�$���G��J��N�(0�t+G@&�+��y�Q�� }����&�^��`-��*�G�yĚ�v�u��a�2S��.���'3@\��V�hA�Wց����f	k�����Aa�_Ab<ߢ�RK�͜be�s���FGj�Z�jtK�.�������I)ʌ������c>	���&�	Z��C�C����C�n#!�-!r�W����F�w���D =(u�A�C"F��ꊁ��!Hoh��1��>,%�4d���,R(C�ØԆ�?=]g��>#��ID�����NRn�׾��z%T6'�1��~��SG&~���D��B�2�u���͚��
���5+�(��}���?v8����E���T��r���7u0�!�u]4�T�M��^L�:�	b�XZL�w	=;J���s�Q'��7�n�F��oU�|��KǑ]C���S���!��(֖���:����5��P���k?�]e��;�nK`��~��<K~y�)md�F҆���+���R��yQc�pa��T��,��?#��Dx�uϙ�V4��;S _$\o�b|E\-��O� X�T����jw�)�rBc">q��Ł\�=50Ucb�%�«H��ݵ�s�؉��iv�v��_٬�A�!(y~s��Pk�8�k��Bm��ب�}/�D�(��"�11� ,'bÅ�KNY��{וز߱�9B.�7.��A6Y�d8��~�w�p���
3���
llZ%�'���b�S�F�}�u�1��x�4pP�lg�]���d����CM�*�G=wG#����D+����Y���3��􏠋1��9L�G�3�	5**��Д�	��n�h���8dus��}^g��E����E�ɵ�����Ղ@�!��ފC���[������aM.���k���z�SRe��s֕�Y�9q^���_���"T��hv��Z�u+�{�4G>���Fg<ߛ��a�ߎ6�FSr�쒌I���ʪ�|B@�3�j�v�bm�p�����o:�뗳�Z��������>�0��iW�?�sOy���g(��$��Xm;9����/,xp��F�p�a0�3-�R%g�i9�����6�*%y�ւ�B]P���7��k���~HfЪ
r��粧R�2(�M�#����D(o�Mٕ�Yv�3�$ �I�a�0/z8cx�cR����'L�ܰ�7D���uvlZ+W�MM�Z��#�C?@��v/o[E�o��Zo񚇯���n��� �=������Н���������sF������r�b��SR��\m��+f�æ�]Cr'Ц��cؔv�f���*g@��7+e����NHEl�
%oL'ͼ?��V�Ҋ��vV�"�`��P��+��M	�E&pY�f<��	P��ߧN��I�<<e�R�Vj%2<��9,"dANŴ�(�綱Z���Z�\@� ��_:���߂؊�(^�aS9e�m��YB
�㰚�w��TK�C��|�a�g�9�j:�\E��]V�G�&q*�v�]� �#���ѿ*Ac6���t/t��}~�@�?�R !���-�g�y�|+Ç!8ŢL�e$J3�>boX��Cr�H]�:�$	nܡ���D��@x�bb�ˡ�9�>��^ ���+ad��p��E����}eQav ��_!;�:������|Vb�*�"����C5~)P�P3�-"TT���2�^���h�T�sj0����|�,=|8�lx��)�Jn��v3j*�����w�$."p�jb���#�O��]�Bav�dX�έuk�6�'��=�9���	>EgX��}G��萀}}�R��~��=��ヹ�`��4ŲGQ�ح�ұe����1��.�
H9�?��&%/��"��K8��U�����1���RP�a@�s�NvyM����L*���O�C@��0��	��;ˎVV�(�,����˾�)F�cszr���� ���_���`���6h��&Z�%�]8�^�G�A�+�Y#^n�[]���[�l\K�p��p��v�oIٯ���"���d>xei�Cu�+(��=<T��v�m�b��=���s��i���E�G���?�I~Ű�a��b����W�	&�����VP[��9oK-|�L��.4O��sg����������-�s��V$�k?#���u	��K1�|�����y�W�Uq<��M�h������
�'d�;ٍv����M>s6������ٰj���	U��yi����n��D����x4Q�"B�2� 8RH��8?5�<��.ш4��;?�9|4�u'޺|� R��b߷����m���<հ�5�O1Y#�(a�`�,B�I�y���~ �.���b�M�*�����\��K��1=6��6|�c�C�i:<HJB^�wiNi�MT؞��T� ���G�y�@veT�u1kؔ0j�7qq��O���h�I�����G����%f} �Р�;���@�D�Iγ9�'b���Q�7r�m��f@�,�a��B#R�&�3�1$ {�w\<z͒Ò�ՂϦ�����Rl�}E�^��;��[