��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVD�6�����;��sD���L�S5H�j.F�0K_[��e�7x��������&�ǝ�+zA��]��~ا@H;�W �v#��s�8��yW��V�>!�/�7��u���nEA�V���E<v��b1Ø^���#K���lӧIA�a�V��R��tv�Τ���i�wJ�'�دv)h�V~�$v�p��"}�v\-8�������>�`)���a��rl�ʩ{�Bf��� ��|4�VDG+�������X".��>��'��E����F�Rm�I�|^�Q�;(1Z �bRw�����IL�+�{Dr[���Ѹ�t�sœ�k�Q�@p%ΙN'�^=79��r���̿9�A�_�@����$�⭜�$�"�T�f�ׇ�[x1@��-{ܐ�Ӊ�-���:B������+]b��)O��<$e|��g2��Y���;��sD���L�S5H�j.F�0K_[��eH�!���Ȗ��h�}D�8����TT	q��$a4�����i�p&�K��~�MUs �c㚂��T
u�/%�ĩ8��[��`�3r�O��C��0��`�R&.1����_0e�v�h�u���;��.~�Gj'$�o��'j���j�r��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���4*�7\��4�/�I����D;���N��j��D���s���ħƿ�9c�1��8�h7H�u�ÍeRuw�C?3d/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�6A�7Oq��{b�2"���Bpш�#w��q�©���B���������'Sea�8���`<4}��(����5�2���[@%����nEA�����G�>�"PT��3n�(�u�����!�M��E�2^Q� �2��m �A?��I\�AkF˯�+)�Ln��S�WT�����Ne�rR6��I��'�Vx�%L���|�r�HzL͊�q���Vǃ���p�m~|�֚?��]t��]|��L�JHn��z�܋�F�]��C%�"�uI��'�h�5,Wlr�r%)cALn��S�WT�����NhΕ���iv�g��gQ�)x�?{���x.�KnqLn��S�W0�T��:hΕ���iv�^�F���.ᬵy����w���BlzL͊�q��1�KB|1<\�5����`Ko����Ȑs(�"�H���o��qo�:��7��k'�w��-�*?�Vz��Y9O8A( ����_�h3��{I���s iG/����׈����Q��K�NI����y�~��ۢ��i��>�`p�m~|�ְN�@�#��I���'��=�4e=��-������yMK�o�Yp�m~|�֚?��]t��1	�<����)��0�E��zL͊�q��UG�s����5����`K��;�R���5���T���n8���ٳ��溂�U~܎VV��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~
_g��c�_�s���H{װ?�p���H�MPq6.JHn��z��p�Sg�3�C�u)�6�Օ��qv��3�.�J�}�|�݌��r��VYW\E�e����KH)D�cn]�#�ڊ<?@Pʶ=����s iG/���������&���$S�ݪ��1#��Z�����XP��ȃ��<2� �zy�g���+�Ȃ�u�.�1�a-���7a
��r�Ln��S�W�'!����è�PA'�(���B����_T���a�aq��n����̞��>�nQ�rV�� e�g����w�K�	�<���BSG�p�P9 �W	́�p�m~|����� �ܰ�a\Y����+���LQ��b9����pP�o�2��m �A?g�{�]4�W/S��8(�E���Kt㲎�������1#��Z�����XP������9�p�m~|�֚?��]t��N�����?2{���zL͊�q���ӫ��%��J����ϟQ��ǺΕ�����a�g()��ikp���H���0H�YS�T��ġ��,_R,T_<�3+p��@n7��k'�w���j����rN�ǁ�f�TJؓ���!��\�v�q�C���z�C�f�����	�vI0���ԏ�.fOe	�Bn'g,��Қp%���(�6o��q��/�����a+Q���f�,{P&l����~��=�����A���ۖ�92���nQ�rVe�Y�gtH�m���E�Y�!|�α+�5����`K��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xS��.j����#���F�e�z`60�F�e�F�Y:(�
�*S�I))����A�m�(};l�-��Ln��S�WT�����N���G����Ћ�l�T�r�&U������G|M�1#��Z�����XP���pZw���ƫ��Y��)�gP���L]&&�@��7�	/-�I4��欱���j���<����&��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�I��Yq������I��RhF�䦓������hY����r�?�o>�3�lrև�"�GI$��ǂcY�~�s<��MR�ɧ�	tc&�j��1�a-���7a
��r��L;Л��|#9������/��&�[�$��X�S�wS& >ht[�����GI$��ǂcY�~�s<��MR�ɧ�	tc&�j��1�a-���7a
��r����~v����"X��[��Q[R�7hY����r�;*�}Ւ�~/�O�	McV�6IWJE�YY���F;�I�e�,��V�jQ��r��#�F˯�+)��L;Л��|#9������/��&l�L��M�,���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8�/ #O�)�+���LQ���"X��[��Q[R�7�=��3��5����`Ke,fi�U�ž�'�t_�GZEh5���'n�^0o�hŁw:����v�8:WsS
��J�	�LÆ�o�P�W�2��m �A?r�ĵz��ݦ\�t!�ǿyXAm�Ln��S�W�כJϾ�ig()��ikp���H����5 Zm"��;���Nv�/T�`��5����`K݁.�q�0��E|�,1#��Z�����XP�����w�K��b�����(`��ү/�O'�=�!|�α+�5����`K<i���A�5�ϟv7�ܥ��2�\Z�ؿH�jGjh�rO-��B'�P������R;��3�lrև�"�GI$��ǂcY�~�s<��MR�ɧ�	tc����1��;-;*�7��;mQ��8���/�6	�4bpP7koеI͢'�����t$I+�V�6IWJE�YY���F;�I�e�,��[�9q�Y�{'%s�h�v��T�v��1����ӯIJ ��`y���]���.�#����1�,��pϓpy%��|�����V��ߝD9�{��灊�O�i��ԩt�t>
x!��I��A2��m �A?��V �-�n�,��v#�[�l\�;���[����|ʘ�{V�K�Nv
wHp�4}�p(��ou�sz#yZ�����n��BI�f�x�4J�P�3��������$��Xo��I;��?�*���T��*Qx�Ԅ��'n�^0o�'vX[��vW4��`��Q��ǺΕHaU$kX�9 �W	́ܚͭ�����^��t�������QOm��/a��\�vŶ�T����+���LQ�x�m���#�	�Zz/pQm�I�~쀨����Ћ�l�T����e!M^С$��JHn��z�F�x�aK�k����k!�M�Z���	���������zռGM�r�
b����2�W\@��u(��}/�1�(�T<��y��j҃�d��ξ���e�J�Pn\��wg�o_����0@ȹWpH7���
I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z���I7��-5r�p =(�a(􆿳��|�vv�po守�u����kL���v��ٙ͛��#�e��H3��i4�0K;V&�٧��;?C^��N~e3Brb��&'�* ��z��K�:��x���{^r�y�����@���ɬc��WN���'nZG�4��K�GI@1��i�װ��E2��m �A?�|����1�Z���=�Ln��S�W�כJϾ�i�I7��-5r����%c��P=@Ч)���;����U�P�0K�*���"�"��|��R��C� �`�����d��oEd�\�-tK�ip�m~|�֚?��]t����nH�W��b9����2�u|���U��+�Xa�H(�˕,+*ͮ[��N5m���z�@ʶ��t�K��L��z�Ĳ*#��5����`KVkLs��dJ�+���LQ��b9���Ȓ��u׿j�h�<��l���ґH���'�~��¨���ې�5��W�/�
-CȔ��Ћ�l�T�Q��O�بeD�I�1#��Z�����XP���#���1���Q��ǺΕ�|7J���UR�J��\�}����� ���U�e�7����	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�����NlU����z~���ӯIJ ��`y�����(��u��5����`K�z~~�Y_"R�W�u+Yi=��o�IÙ=�H�R���}��M�+��l~�U�{}��*���M!󂋷�(����C4'n��=?���͞��>(�J52��m �A?���"��|���it	�TU����z~+Yi=��o�IÙ=�HVkLs��dJ�+���LQ�{p�uR�R�W�u���_�)�Yp�m~|�֙X�D��H�MPq6.JHn��z�%�,��CU���it	�TU����z~����.`Ϊ�/-T)x�?{���x.�Knq�w�'��I��'���h;e��w�5�ϟv7�ܥ��2��&������7�0� ���������n�T�?��4��y�-Ղ��hV��6ۿ��K��a'T���W�J'�s��4b�s��<�6�Q=Zʓ�p�i�i��О	Q��J/[�M����`H�ʤ�ܔn��aK7��������ђ1��{��dP��a�Š��7�"��r%#W1�Z���=�Ln��S�W�bOM�P�CC�`�/�t�+y��y�$��Xo���f�xO�Π��yGb���n8���ٽ��j�Q%��{S'����x�]?q�����f-����0��V�6IWJE�r���秹�3I^�v�[�9q��q���U�|L�P�i.��Y��¤լq��/�NI����&�ߝ��e�4�+/r��bQK��Ņĕ|G���r�����+�va��2鍔�	g\A�Q�Q&��0��*y~��5����`K-�U�a�&3�W4 X==%�4Gne͉�Xk����0������Vϓ�;Zr�î�D��WZ�M��x�	6`�Lլ�w��������.�学u �$��Xo�J[��K���2�$����*� �d�Q���n��̒��b�|���{�\y�.�^�h��Mޢ\g�������1����r�x,r��0UwpB������õ���:�v���)L��mU�.���[;Y�@��O���Қp%�&zΙ�[؆��Sw����Y%�����n�uw��z��v� ���Y6��&q�oldW�pv)2O!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(]:�z������+�̣��ަq0��
�k�� ���4�Mޢ\gȟ&��s퀹-�[��y!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3� Q_dʥ����[�H>�ɨ�m���y��V�	,���_s<��H�;� ��kׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���A���Ձ9�N�c����7�}����)��Rbk6kR4R*��Ǳ`��W�gǼ�\v��؄aX܇5����`K�������[�Zl<sPQr�2U=e͉�Xk����0����AH=�3"�q~t ���ue���+>X�M\L�">w�"#6>^�`���U�`8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��tn���x�Un��]p�}��ī�v��`�7�p(u!�^�YH��SaJ��IL&L�8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���?p��*-��M�B��GVDs�i|�)1�A�7f9Wc�^}�O7,�m���.�D_*y !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�{wx�m^Br�hM+���XC|L(�Nq�l�KE;J�[ҕ���*�Ǻhu/
e�Q�o����CÏ'2۶��wc��du˷
���S�|�Ĕ�*x�j>��i6�0w�mL(��ߠ��v%�T����1�2� D �����&p���7 O��D|��ϳ�����i"���I��'�;���6�?|��ͱ�/f�6's�cbp��'$��O�&��o����7ڮuK�i�O�ߖ tm�:�'2۶��wc��du˷
���S��ݢ���j>��i6�0w�mL(��ߠ��v%�T����1�2� D �����&p���7 O��D|��ϳ�����i"���I��'�;���6�?�ا�	��/f�6's�cbp��'$��O�&��o����7ڮuK�i�O�ߖ tm�:�'2۶��wc��du˷
���S��'���1�j>��i6�0w�mL(��ߠ��v%�T����1�2� D �����&p���7 O��D|��ϳ�����i"���I��'�6���ퟓ����e��47w|s���0�$i��k��L[����Eۨ?o᭹�A`9���^"�}�g��a`ծЖX�+/7��xƯ�)tP(���5��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3?�dq��U�f������K���_��"!?�W Vo+5K� }�ħ�nE�08X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�FL���/��p}�6�r�Ա�J&���w3�#�T�����y<��I;�ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(]:�z�~����(^b�㷊��B��h�M�>NQ�q�l�.iA�$��Xo�k�Ԧhg���E��Y���N�*}*�@��O���Қp%����uO鉧xL¶���%dH���[�G�;��:P��~�{��P�ڇ�U3�3�����Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��� �w���teλ��<�{7�'BWG���a�s��4.va�M|uŒl���F�sȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3	���P8����G���Ģ�?Ex���n�Tco�������V��jڋ���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�:�rCl �����&p���7 O��D|��ϳ����j���