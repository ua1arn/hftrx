��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y��� mQ{��0k�Ƥ�I�x�ݬ��|�>��'{����YgBK�K��!c]�@I�2�`�p�`��m�M�L�f$�AJ��KM�,��x*������(d�|��F��6�\38����CL���3J���@�z�ʴ��G��/	Uы��|��{;����,[�@�Y'+Z� �s�m����+;J���TNͩg�e��`H�4��߳����U�L� �s����qVi%��>�2����[�X�k���Pv΂����VT�;'B�hQ�o�����/&o�9�����A�6>�Pt��(�O3�Rx���?^���!��/���Ko�W�c^�s�O^�C�r�,��+ؖ��ҽ��ֆ���h�:�q�]P٥��t,ݻ��3Iq���@g��5&�l�K��όL�"ǕE�0y��>�[������:�M5%�V*%Z�O
�ܘ�>E'/	�u��-�}��v04�Ef��L�cjU��)�9�u=
HD�1w��@f�1��yy5dŒ���B�y�.w��G��Ĳ{y�x\vc!�+-lf��d@����aw��Cֆ~D�������~şCk�4A��9��B�*�x'�����W[@ۛpe/#* ����G�1t����ɇó~�u���o�o�����Z�)c�ݏ� B���3�|,��d5?���$<��:5�g�^7���7�~�psj=��pP��=�lz-k�X2�m�� �ĂA}���.���o�R]�5æ�^�;b�?���^�/*��� ��
��ߴq��Ű���M�)?�X~�<J�SA����/����tx���zU�K�H�;�'@�ek憋=��������QK�HU��+dؕ��H���u�Şt�z��'y)��Ġ%<�dc��{������NE`e������� ��W�� ���v�{B�Bv�!=*����Ο�-�F��q׹Z��\�b��A��8�g������#N½_g���;�R��f�#p���P�H��m���2$AHc-fδ��������A�@@��\n��<߭s��>2�F�_&����@�Snap	��.J�F}5��w�,К�-@�o��� ����<� |P#��^�#���sE��	B��&�/sT�69�S�M�_�Jq��	���&��� A��̸�/�N�yJ?������O.�[8�@vٵo�?C������vCD��[�Z5�u�0�P��s�NC��I����c�tiTE�tK.�^�Lj-�E�㱼OU�_ge�}������<�U@X4(n9� 9�����&:��fR��$d�v%���:���-Ν:��rWH"Tp޸�s#��<cG�	�I�9�pd�[h���*p��2 NC_�{)E��
,�{��#$�+q�X����$���b���Jd�=4�
��������.���������]���@6�C��̈́�/K�r��5.�C���N��N���q����_�!�ONdln�,�����mK�A��� ��S�/ ���CrC<�9��������e��Ӂ�9}G˟xӎ�u6
Tԋ(f\��C�F$�gS�٬�:zW\썺�9cܧB�`���(V;ů��_�S�NK�R����aq��W2"/Z�����t	Q�s��x�L��
.Ծ�M.�L��)+U
��"h���qf%��8�+��|j���ORl�&��pv�L2�yL��u�I�a_�]�Y��E�?U>�=������%`��Sl�C�>Ԏ�W�j��u��W��Tp�:t�f	5 kc�%�sD��	x��D�z��r��^F3�6�}V4X���z��Mܔ�g���j:��&�=�
+�$Ee7�Yg�?��E�d�o��T)#,}~[��)��h�	�(@4G��Ձ#�6|YX��;&�ߧ_��&�I�J��|p������ԡv�������<���*-�.k1Ӿ����b�i���M$-������F�T[�
B�Z�{����e9����(ڞR]�I&{�C�主���\1�i������&���1q~����I� �'�	JD�C�{�~媶L��?&���3����Vu��m�V�z2ƻX@�N��-�����׹��M��wg ԇ�tʒ��Zhr!vcB�Gl��N���,COޔޔ�E�P.��͜�*n=p�ui*+pS7gl-��kr���^'�� V�f&\0���^�x�d�!Z$��@���N��s��<z����H�=�x��A�$ݓ3J-��ZL`��Q�U;W}>��#-k�Ϭr6��U��>�3�,���{�+�ho�O�5B0��3���%b���w�^dګlܥ��P+��x���I2RU*����!�_D�����۶�Qu�8�V��ځ��.�U��Ԝ��Ѯ6��tY��:��̻�y,������5B�v����>>��5�U<Z|1��IDY�~����O�Ya7����� UnA듏���$��+�)��6Z��V��-[RX?=��&�����c�s?z�9l~튐���'�H':��th����*�T؎e�A\�!���������Ro�*>	���*����s6��'b�Zl�Q��4	���jD~���_�ݭh�b��m�ZY!�R���b�p6U���'��#�E�o۝TO ���y.c�~����7�=�
