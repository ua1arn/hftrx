��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P}*����]�/�Ϗ���{����p���ȁ���r�C��9k<����Q�ܨ�C���t�h�������Pk��=M�^_�:7 �L�����$#o7l���5�㫢}�lhM�#Ĝ�zH����*��T��C�#d	���f�^�2�����;�(����Ekxb?ߎwg�k������t��{O#D�����~N/ȷ������Q������ �R����F0`�FF)M5}fB���a\����0"9��}������U��9�s���Ajq������F7f�P3?�X�ê l�ٓ���Ҿ�I��� �w�mG�,�(�d\8�N�Lh_#�7��RBeTI���wb��ja:�#�[�@;'���`��z��wa�F��tiD�vG�Tm��g�}��瓑�,��[�|�^h�q�������~��ڰw;sS|�
KHԬ{�D��eG����j���J%&�7��?�����I�K�Q��Hl�LpC���;��91��Y�AXE��ȦF뼝B�g΅MΫL�h�@m�W���Qg��g�Yj��[���>a�'�b!�k�ڂ#Pr��W�$A2iz���h"��oE���D��% �Oa�a8@��WO����B��ֲN)['Ɇ릺)f�^>8���ի(�X�)���D�P/�*�r5�@MM���e�Q+��F�l���] ���P�}b�t̵���\A@���Q^���!3��'*.6<-7,��>欌���;M������j�a�9��L�xĶ�z���,u��  �A��T�����5w]Ԭ@;�b=r����~��%1ɰn]E��1�N�<�����$��i����OCʦ���8�k���3�� *Ӫ��I���\�D�Z�S�'l��^�S{�$q+1k�R#�_��v�C�.8���|38�m���}�}t��܊��]^X����1��e�;z$���g�s�pX��e^��O���p��t%MVb��pl�����=�.Y��ۖ�M��CZ��@W9��-�3�0晽��!{�"�P�~�؉��&I�_�T,�Ҝqf��'`�"��4����FJ�AI@aeV�T�P[8 ���~������]�����je��1g�h�^H>B���s�5�^�,��!���mr�%�@�O��x� ����]$·�7M�bK�^������[� �>t���kj�c���D'FW�MX�Jv2�Ɉ�(�ejt��\�a��}fc������3T�>_@S�/Vag*�"l��u~X����ntO��%���G����M��z����z��I��5g�b�s�����u�,ht(�yEv�0�2��M�<c~q��z!�Y��9n v$I(������j�{2�x�6����tv�]Mo��:�+Arkx��M�@�,Ca��K~aV�]GI}	Ӕ	p{�+B�dC�J���r�� ���؋�cm�oL* ��U?)�Ø�I�I�m���;����O&L����U�S��f�u(� ���R�8��o�!��Y�8t��N�G"�mf�{�j�,�q1	����h��F1mWV|Q�H�3j�)u�L�寸�〺�L��_~<���..�'��D��jR�[������P�Ոy�bB��:�6��i[�mr�]�J�Q<���oU�@?H�̗�2n�
�C%�������qb(����	a7�^2����* �2�L3�
U&v�9� jwk|}�A���NWBJI��pq�c�%/ݔ#���[��*pDIӱdફ�ÿamB�;Ȗ@�I��zc���Hb]�c�����Y�m�K�ғ;P	�j+��l��m��r>�1#��Z�����`�b��}��)g����;yh��.&� ����0�~�<�(��۲��5�p��r��X�)3�����J�n�ue)PoN�Qk�v�fm� ��qoU|5r�_���[ހG�$wx\�y�U��(;E_�{V���\��i��<�FE� ��o8w�M��e_[Q���Bx�~� 0�zV���d˺�ѕ�yS�Z*p��,ke�A���mRm#<���♎�#����@�#Yh~� *�K�@�jQ���M�G�՗��D�8��$�3g֓äP�Y%�|�,hEZ�� �
(N�|{�Ú�W�̊Z.+֐+��Y�J�@�u04�oE �����Q�L��c�rM܎6P�EN?\'[��o{'����<H/�s�s�=*1�mP�ݞ��t�\��O�����'.�_i4�]m��W'9X<�����X��>-	�x��6��Wv��tmS���O�#���p��%���_�}@ �MP#��g���sE�j��'�e���HY{���M��1?�.ۚ�Kﭪè}�bR�(s�;�e�$�'�LAeܷ:D�Jv���� ��X!�_�ϩ�m"�/��;�} C��A��TP�$C`�%�("��,]缤}Q��-:�s*�U{b�������+���:��z�PX*�4��V=���\U��_'S ���u���C����(2���us+��o A 8YĈ��[�H_A��1�_OHi�T��VM�����H�N��\�<�����t�h3% �-G�W��R��ʞI%gV̶���;�����'ē�*�V���[Tbfg9V�-�W���m����*a����ح(��ņvWe�^YA�uK<x��gB�=f��x��d	"1��k��2�On�rq3w�����y��䔱g8C�P���C��b|�Yb�~<��~�b�\���h>���+�DQ��uт~PYF�B!w�@�<.yN��L|)��>3�y���є���K]���uSP�(��CV�w��e?pJ��G�����j�(����������9�z��D
n8N���m��mi�����|�B}��I%�$th���I[&˥�bJ,�_X'�ן2LZ:9)�Af!�K�,�N�5�4z��T�aI�cb� :���tUmb�9B�c�'�"�;(+�V���}d�
2+t��	Κ�함�n2*�>�{�;�DM��/�~�H�|�rę_�,�G͇�Gی[��^/T��Y�n}H��1e+7�(�D����q��Cu�HJ�yweb��$>�r����
%d�BJ
�뼌i����;�_�ge��.��.k;�Y���|�c�oִ�oE���4`�ZW�腥"�5�-"���!�- ث��9(Z�}�3�D-�L �����������	����~2�%3fqrI��]�aZ��Q�NN�4*��vydW�T)��!d����dj;)�[?�v��5;>�C�Mz�m�������-�|�to��B�ð��	Ͻܾ;�YG{�����9ԬС�窯b��ní�8�[<+x���߬�ab����q�*��@�7^S���ϾOO�;�]����&�cU����������yPP]1�NU����Ua�)���N�
ꖟsγ�eQ�H	X�_� �Y��+��G�8�̕��`��k�kQ�W{��?f_ż?�����9��v��U����˯}E9�$���ѕ������xT�)�>������H��)\�����믡��n�U΋T٩��yM{j����藗�}�u}yX�Gul�,������Ob� )�~���s��F�d�{ջin|Ln>�fX��A��3��v	�rZq�E2W@��R�Jr����^�ۧ�1H��S�M���`�Y�;�ܶ�/�U�Ag�Ѭ
��LM\���eW\�'�%5�<��h 2d���=���i�0�,���O���dUWL�ʅ]dT)���(����q��������,�,�!�72��n�`n�/�LfE4�Vm�}�h)F}O��qx�L����/�Ag�v���7x���S��m�pё�/(�j����ӃȰ���V	�R�5�}�u��9jf�����(��O��g��� H�+�*�`��1��U?+����i���k@.\�5�y��O`:+�I�����Gj��. v��Q��7hD)百C8Ҝ�<��4$��@N�	�-{�]�b9L�/P��8y�(Y�g^Aۥs��ǟg_(��/̌|��,J�4U�T��zL�����1� %�R�f8��~�2��������W���FwI_{�b�򔪩���I��ֿ-t�nO�!w�޻�t�o����u�z��o�WVe-M�0d}$h������Iءj�눵��{}�.��J{�4�8�꣐ה���A�H���?�XS}l-��'5����z��*Em,x�$FB�H�M�l�"Pw-F6��h-�ΐe�s�"�a�VO;g�캾>Ȥ�H����qI�#������LS�b��فu������T���Ѩ�]%Q��4��_���6�S�FhJ/��_(��i��h����//�T������S�E@�}���?_���71��%�ldMj�u=ʿ�6�w
��t�h����IӟM!���C1:�ˬ2������q�i(��|�����C��v��nHU��hS>r�Z>�<O�_��D?������Zs2��{����]R��f)~U_��L7�QG��хո9Tq���k�8�m����l%!���7ge�e����;��m���Ɛ�[���VS0���)�@a�<@�e�D�ׁSD�>�:�\En9���<b�����ɋ�Q�oJPdcPp���P8�hwa~s�Ըfo�.�Q;2�f���y�>����Ֆ��$����4gk� ����vН�Z�s������*C0L�QJ�p�	���9 ����\�)�?w��E��#S�wr�����]���ă�}5D�}�X@�{U^��`g�D�ȉ<L���3k�ޑr�)7�櫭�2���;��T9�o��3{Х!�ځڞEg�/��k���#��0��g2h�W�X���X&V���>�p<�Q�Nw{�9��-F�*�H3�Y=F�\6��f��s����kF�kJ6[��:����Yb�s?7�5� R�O����$��y)u,� �n�ٞD�Y���,�'�VR-���r��z���ң���{�Ar\�'�	A$��� ⹦�4 z��">�J��9��Fo:Xu��:��X�f#H�R��R�&Gt`ތ�hsw�\����eūf?P�x)K^a�׏X���eӽ�a���Ł6nj��r�B�G�&}D�/8�}���e`a�i�hR���7�{5h|�ѓ��&Ҳ?��-'V�����N�PS�I���V ;3�~< iǊ��b{�7u�~^A���tBA��z�7;���V�B~�������9�0/"���gDѮ7�[�������K��l�	��j�m��1�G|������ڿ����}��=�6��RI���tX獘^�w��"s�����'����L�h!v�('�F��uOY4,�
�����izQ��{;:�iQz�F`
��,u����|ݶ'_�G��,�O�|�k��a�AHL�Ʈ�M��N�n�-2 qz�7��E�zu��?[	�H�D>�-�T���D�^�B����${��v�(����v�.�ևV�e���O�	�,���p~1�6�bCv%�����ޛ�>_�(�q-�	. �Uw�]D6֚W��	��9�rGjm嶍�\8���
G싾�[P��Z�߉g�b؃�~'��{��B��mU'��4���vU��s�������SzR��/��i�V����W��ݝ �I cb��P(Z�� ���Nٜ���'?�J=�V��4��,�q[�m�I����Z%���o�R�N �/��}ޯ��� ��֜�O����a�����ȅ���	��F���6���س����9~Uq�x�G$nם_�P�����eL�2��E~�������#D8i�� ��m��:dj���V�x��tv�S����	�T�f���A;� *4M������Z�'ێ�)� ��wÊ�b��."�*+gp��n�v�o��Pf��9�Y-98�'=%��0�l0��/bF��:�0�d ��"�w�^�)���Ozg�rIc���4�Mݍ���J
-U_��A��F�����eN�厚�es�k�\��~��ą6�^�6���v���U��n�M������a�c�n^�I��R!�����0ٻ����	��jA��ɉ���F�E��9�mw3�mUJ�j!�̆�%	��,�h���F���'K
�����Α�3(]�yō�Rv#I��w�	�z=/p��-Q�D��IVVX�������
�i�Y�a���ۨG��DWjl?�}}���nEQ���.V��p�eLd$��Y�Ҙ+v�Q��aX��S��>f�n�e�fa
N��^�h�Oռ�v����N8��q6��'Ϧ��qG�1jN�;I	'�$��<_�!���������r��WA�N3�v���$��Z�!0����w18]"qw���A��+�a��$5;��~�w�m��I� ����%��Z��r�Ƞ�"����˧��gȸ�"��ݨL�]�����;��۾x]�x��c
@%�lc���m�N�����	�sRo��/9V����^k�|l��U��X�5�M�i�P��Z��a��a,!��qh��Z����d��#xF��e ��k���H��'�-�k2�h��_�H�ڄy�����h��P��3T� �<®+b3t�D�N&i��S��,a?�O�8�5�.&�ꆐ�j��٭H=>!��h,�įnT�=7G��&�I�N��иkW�����őp?��g}���!�p%ՔÀ���V��m�Ɇ3@Ƌ&أ*l�+@�����s���:�2U<K���?"*�z5׎2�Ъ(���u�3��վ/��*��5���v2�o)����5���]\�5xP���[�퀽˵7�w���~�Å��o��V�P&�U�Pk�^��!p����k$�1��x�@�@�#�п�7�?�9ҁ�ָ#�ԙ�x�Ԛ��o�	��o�ȻG��X$�KS��U�7��OCyE�3���R�/@�Vp�e����Έ.o")�a��cMuߋH��n�J9P�[D�Gi���گ�<[�V�H,	��?dQt\q���x��� �_"����6j��g��:E��{�����p!Dw#�90�I�v�7Ln<�N%�'/��'�M$��Є}T 0F��
'��c�/�k$Y���sX���m�5���nZ'ѵ�G�)�3>`�%0�O�^��D��H��X}[a��~}��^B�-����^,WՌ�[I�}�֏i�N��Nm�S�u��R��/�,�V�
%D��X���r)Ad��~�u��@����U�Ji�x�"��*�|��-Dq	���R
�8
H�ti�	2��+�P?���q��Z
v�В��r��0���*�s�� ξA]��L'Ay�$Hd��E��#�xV�t�eN�m74�b�cj�U�]�K���F(AQ�����dg8���fʲj�s��QV4��C� N�K|��÷��D������N+�9,oZゾ��{��kCm�5��i�ۼrW�p�q�ݛ���Dم9f����
��F�jC���W�K;� �x��d��tp�����Y�����}��p��q��z���+������@����mh�����
�\Q�����������X�����-ٕ�� (�����	Z�k�^E�ܖ�|R�E�0V����"�����#���z�L���5�qt}6�d��{T'=I�N�,���@�#�93�8̻{���0��>"��;m�����!���f�N�u����at�if�֠X�y�6�`�Ulz<)mPvm�S`�2T���Q�}�b�%�M�n�{��I7��H�R��Ю^�%�yl(:!f����WSA��R&BHt����\���~�4��x�K�o*�@�;n�%�ƹ.��~�+23�����%P�Y�/�-��ոy�'�b#��q���jA�a�-�Rȇ�2���hJ����*���z��^�Ҿ��@62��UvƖB{�����J΍�nF������
���%4h$��;5���O4�ǧľ���yr���X8��l�9���p#�t�V���Z�j�!��pþQQ��IQ���1��tߩm����P��m��j��g+짢������AI�k��@\�DLs+�`f�;*�Z��@�j��E�*E���a�r�_�]�kW��y�a��	������j���]�to,c�P
�t�mQ{�����/��ဵ����ŉ�)�'����\�Bp�b�[�m�C�����s��#��{��Y̲B��C��)�qk��Rt S2�O����l<>)|[��Ŗ7��+�$�0p�>C�R;U}p�&�����n��=�B3u}lR���%�&���~A��0t��`��������۷8�^S5���M�ߊ[�*3�FQ[�8�X'"1�3��c��c��=s�߀�zD��.F?KNWX�d��V�T ���9�6C���:������p,�[,Ĩ<�9��h}�*-q�~�6u_^d�N�4���>a���D>J�w=��6��$���ۤοnw90�Y4�.�+A?��c	U������Hvh��{��(�
h
��Ba����RV�V��4a���5�UJ@V�ꀾ�<L?�Q`V����d@ �o6�����8a%��P�z�����/�*�Jv\���a�xJWlQ�XQ4��u�~�{��������#ؿ� ���h����`rpT����	^��C��D%��0}�����Qz�E��4�w8g�U��[=�)7�b.��>���p�Hl��a��3�~5S ��؄��L|�MꦯEN.��S�
&
�#��!�_M�rE#�\���:�
�
�㔖qI3�3�;�>f���.�($rK����R!��a 7�K�-������f9~fh�%����xKr7�x�M�+�F�0E.8z�UZ(�����b$�Y#>e�+�M���5��(�t�~��^t:����<Z�4�����G������0�y)�^�(�5�G�L����}�0y��Z{&�o+I�l��"�?֟�R����>1I�[�p<�>@rsׁ��w���%W"S���%9hNn�$v�,3�u�R��[���V7�^M�`�&���	O?!�}�-#��a����3��
��T5"Zu�P�3o��ݿ�K�f�dC��i�c���@���0�0P"���1���n���?
x��~ְ��H���fɻ�����;��V��u�h������Z^�rk�W�X�>�[I��K!�'5�y�gt��#�v��'�R�����~~�����͍ݷ�l@��3�/���r}e���ӜW�;b�f�N���6���{S��<����?�A�%��*"�/{N�Ŏ.�mZ!<����԰f�-�<"��ޡ����1�����Ev��*b����k�0Ut�|Vs�����,�t�T�5���e�U�g�8i��e�"�W���ԝy���U�D�o	߾D�;;�G�F��>m��q���%8%T�1T(���2$��|nx͉��h~Sm��<��!��o�u4>�쏂��&b<�W��	��N��+���}�����~��N �2�Q4(�}�DZ%�Ec�V���'Z}7��ţ���Kܙ�G���l��Ȍ���ߠ7|	��Le*�8� ��Fk_�X��**z������rk��x���H9D�7���nr����~ֻ0Z���Q�D���;O�42�����}Yj�F�ӽD�x�]�m��xA�F���+_zP�OTZ�%�i���*��6� �{B�[ I�f��G�}�:p�O΂��C4�¯鯬��e.�J���+��6a������������m
�K4���o��!�.Q�;-�x*��f�'�S�����zn���i�n-bNH��1��)p)��ň�4 ����2< ����K-�1ă��#�l�BG�e���`��z��z�\��Řh���n�`���6]���f~4�4Ӡ�Y�Bc?��!�t�iH��9x��+C�Ԋ������982�(��J�ĕ|���m�y�W�u^o���(Qd@�5����|c�?�hm\�&�(P�����[i�c�H&�fR�����;�rǓ{���L���m-�Dxy-'K��P$��v<�O�GA���/�q)�"s���iXvV�hZ�3� �$lL��i�=oj8����0�p}ow�[���Z�'����w'�.};�	�o������[�n"��n�i���2GÎ�+!����$MU	!�N'�jmc���ZK^��}+�m����yG��T�Jb4y0��Y�ׯr�V��3s�Зz��$���P�X���!�0xB2ᗴ���!��ݱ�S��\Ǉ��U��G�E�˟bW;��O@�Ny�m�k�dHɚ�t�i�2�)��lӵ7㠼)v��RH c��T��Q�
�bT+�#�W�]�~��s�a��u	B�⻢':-���utakN�Mò�Mn�"��� ��c%�u�U�|��)����r��1S� p�"=��R���N�,r/����[z���+�7�x��!a!�j,$;�!h�m�R�dY���7�$�C��v!ħ�މ�%�2G���TC�MI3�+*�s��+��oD��7�ݞ�:G������M�Ӕ��p-����1g[�-��@13M��8V�]sݠ]sk�/.T�A��7ٜ��'�ΉT{��|+k���$���g��8�x�Ň���+�o+�Ǹ<|�&�O�tNP��6��3�0%���h�xE�a�9�Y!a�v�+�_�H�L����o��,t᪂ɖ�f�����@�w���	_E��:�����Bb�0�%���Gz�Yj�S�9�$��zyQW�m��4)���)��˷��!Zz!���%�����"Mo�%>`�,Ͳ�|��b3t���#H��.����o�zq�XF�'��\��VW�M��A�@�5G�l�[��l�d��9��
�ѐ-#����粼�!ހZ����gN��UF���HN<j�9`�V��KZ�E���ݒ�9��-�-q����a�����0	㞻�BO�Y�������?g]
(�8wjhƥ��ez�� ��P��4̗�/9�9TqQ�y��JՅ��x6��Ea���1\�������p�c.�>S#��]��w>΂~��\�I�� iG��`��VI�UrM7������{-�@�#�����tQ�Y�f���K��tƤvv�G��jVi�_רE,�j8�3:���؅�6��6���=��Kd�1�tP��5ؑ⮟�Bq2�n�0��ke/} �`W �o�H�k�����c�8�8Q�2�}MX{}��F_( XCh�~]��� ����?^��J�iFVan��ZZ��!�f������K�X�/�9� �=��vF�iU`�X����kPU9��@l�;�� Rˤ�cD���M5����spn}�d~,�>{A6�a�"���Ô�5ᐲ�W*��2_�|<D��ӗUo����5��}\��²`�����	j�d>���kaQ�hTC'� �;~3*>#�k(��p���u=�HS8X�˙SDS�C�w��<6'�r�[zLY�����1���8�Mg��So�}����w��ϗ���p����T��џ�`�u,L�)�h�}���˚|��w?h���t�s	Jwdt����6<|3�|� PV�Fl{����) ŗ�����Z�ַe	BeU�W�>����0o϶�ca�ok� ���Í �T�Α�>�/���}V@}H�͸�+���B�c���Q;�I�^KZ���rX�'�x~j}�s"��q�Պ#��ΑN$0���
��Z�Z.��ּ�o�!+*ye~���2������ x]���sx������A%�FP�[�Q��2ǽ�01^O~h$6��dh��b�0�/�N����Z�<�dVp���W#���� ��3����B�<b%`g��)=�-���:L���*�"ZR@�z ^j���#뢅u�-����ͥx�U*O�.�bB[
�����#׹[f'����#�W�Li�}'ַ#�$����f&�ŵp�h􇵕�0=wE\
�E��l�gd�<F{���K�8��d��&(�����$��lkFQ�}��o܂2x%��E�:Rv�pb��<b��r�G$�/�������e�{�W�P�hv�A;O�q|��1lx�&�/\��?w�+�I�=a���'�&��W� "uY���<)��z%��r���5�!DR|JOF��{tYJ���zhٟj{��d�z���"Ӄ�J5��)�uk��ـ½:��ht�CY�f)zm���?��q��q�G�k�*��q���ߍ��5�,�Ęʔj�]�/L\n�/�A������Q�0�I���)�������I=.�s,o��m_�+x�~�/m
"�O1)V�z*�� ����-~wuxE�] ���8N3i�N��3��IRjY��GQ'ڽ�R��|B�א|��a����qz"�%0�x��\R��Hf�����A��њt���;�Z�&�=U�ƌȔ���.Pڑ<޶���`v��A[/�;���>y�ue�nY� �m��