��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ�E|�$�c���~��K����`-*�Z"�3�ג4�J|^��k��R�b5�huͮ�*r�q���U$��X����WB�+�	@��%�M+��54����j�V���u����a5m"��G���Ac�B��.��Ȍ�z���yAu�Ф�nzP��vp�tzz���\s���H���g-.��>?�sY]ft�)30@�q�!��_gY��.A�'=�v�SP\��z��Q�T���i�:�5�T��nE韞��ξ�,끚�6�����*P\l��#�z��0'�|�?�M��6��6Z�M�+���q�D��A�6�x�e��y��a`��v������}��<Ԫ4��;R��o�	���PEzO|����tzfҭR�~�V>D=D�z�4c�C��G�n��L�7+�QkN��3���(����d��ic;��CU��1�Caţ��p�_�9���jg���}@�?8��,����s�e����/�^������X�6bceN��{a�,/�D��7Mf!N��V"�G�[�?a�?��N:��iD؏�ˮ�$�p�.��* B����G�Tk��+}j�.{�a~WwP���Ѩ���q�VY^�^m	���>w65�"0�2���2�M@6���_(lwZ}�_�x��N�e;���B�J<n��d!	��^�.\X���|(10�+
��5v�Û������i�$[��>OC B�����U	0D�XP.w�x� ��%���G�K##%,�1��-��K�^�?�'$�jU�3DmU��D�/9T$Z"�����D����S�d[�|�.t6K��:�h�q0
��	�S��Pe..��+!�9:v���T����,��0�v��P1�M~èk�\�T�^u�򪋆fV� %Un=�2B��� _\��N̽��������:��@��b�)�K*��lG���F��8X��Yi��m���F%��V:�W=G�Y�Y4��n�7�l/|�x��z�l��S���3�P�Lb%{K3�{ӧ���%[H��@�`��s�7��+���颗�NA2�:�Ji���Ɩ��0uōl�?g�_ 9?�*{+�05�=wŒ�����b����寧�_Z��S���6����Uzhؾ�M*%GPsS�M��@�@�YF-M���/��=(����{^�#t����z���ֳt�<���*�<Ӗ���r���Q`-�5�}��*�H��ż5ԱN_z	�R��k���Q�Y� ]r�͈ӏ�{���m��Z�9�e�LG�7(	��>�h���c&Ct<��~j��iXI�26u�A��h�o�֋2�6h�3�(�$�,т���rD���CLu/��y��� �3��Z�P�C�ݱ�&~TęW[;E��Pmzi'l�]�+���P�P�;�Q:VS�W፰�vs�D����RĹ �-�r ��X��(��$����f��`�W@j��:�gۦAɡ���I+��u4�"���=��? K��ZI_޶_��p3���aN�{v"#>�N%�&�jDg�':y9̬]H�T�PD�XY��"��e����%J����Խ��Z���N&��i�<�y��K�gg����=[.��"6`)������~_�������Dt?�h�x�wyJ�r-��l]�Rs�3�������
�DeN�Dr��V����$��	57�T��{`�X�>)�m�?�ޚm���X/(@��t҆y��D3��;���tF��c̑�^w�ur(S�QRJ����Sk��>VL���������0�k%�p֧
x��mzҚY|�3=T4�G��q�A����s�	���9���>�.��������w���[�,9����@ے`�1y�Ss���T����Y�,~2�G�0��8���纪[���/n^^�{Aoe��kg��a�Z�HyD��[	C(�E*hr�!.�{P!;_�؍��b��Ż�e��ۿX7�FLu5���Ǹv���n`p���bR�5b|h%�)OjB~��ä�7q�&gv��.0��}5Dk����j�C��P�;Ӯy)
 ��/��o�i��h�b"�\W�d*x3;����A��Ϩ���Է�X�L��"���F�U:���fT�8.�U<�R��q7t��%�~{�T�'����Z��'�W�5���1V��Jf*\	f�!�l�l��-�÷5���*�Ը�|[b�P��l��9���!3��1����Gu7쒭z���[�1rN1u���~�s���fOׯ��q4]�,u��,:̞0NJ��� �m�M�áˡ�wsc���kR��ǎX}J��ְǪ���\9�p�#� �K���@�UrZ�
V��i:�ұ3��<��o�k�0e �S����q���LLfD�*Ғy���%D'�
΂/��Bd̑�w@�l:'c�B,ݰ�5�T5���)&����댘ҧ4�)� �X��bD�Z�*��DZݫ�����}� ��#g=��a����)uv����荄�X�w����6�֚':o����<�4n{��G���;�G�Q�a(�c�
}Q S�v��&
�+��t���%�П�y������_<�ۼ>�?��H���T��&R�?��<[	l>2�4hh��.�^R��L��*��l���ǻ/o��x�#k3�"���rZ�}o�cUo��X�Qތm���|�� �0����)���)g�-�+
<Qѹ�`�ʌ B�"��%v l�VK˔q>5n~{Vze"���">�.;NQ�r)����{��4�P��ͯO��
���8庫�_B�}����ˍОP |�F̆���hRBk���\����F�a�1�������	X�I�_�z�n�m�H��D�t����}������إ��T0���g���"笄�{=���2�\0���P�AH�\ǭ����,?��Uu��¸G�խ`��i���We	φ�T�G
���AŤ��Qr]h)�b��̆��B����?N���lP$�g��i2�}��G�����>b�n
hڐ���́خ(�)�T�2T�%�[K-9�^o���APՋ
����-v>)���/�\�qy]X�|d�p���։�68e�?N�уŻi�����!@1�w�Yɪ����_��`+����Y��VP�!��q��M��H��W5%<�9�!!X�a���$ߩ��;�0� ^�eZI�z���t���;�H��[vw�S�"���� sß��(1�u����e��Ƨ��
}�!]�IJ�C��3���C��aG.%Ho�0U�6~߬g(�G�^��K�9�q��� *�G8�1��5�m�g R��6�`��k�m��b-�C�`��;�����g�v�"rYP��)@�����Łi�Z�]��