-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_out 

-- ============================================================
-- File Name: dacout14.vhd
-- Megafunction Name(s):
-- 			altiobuf_out
--
-- Simulation Library Files(s):
-- 			cycloneive
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altiobuf_out CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" ENABLE_BUS_HOLD="FALSE" LEFT_SHIFT_SERIES_TERMINATION_CONTROL="FALSE" NUMBER_OF_CHANNELS=14 OPEN_DRAIN_OUTPUT="FALSE" PSEUDO_DIFFERENTIAL_MODE="FALSE" USE_DIFFERENTIAL_MODE="FALSE" USE_OE="FALSE" USE_TERMINATION_CONTROL="FALSE" datain dataout
--VERSION_BEGIN 13.1 cbx_altiobuf_out 2014:03:12:18:15:29:SJ cbx_mgl 2014:03:12:18:25:18:SJ cbx_stratixiii 2014:03:12:18:15:32:SJ cbx_stratixv 2014:03:12:18:15:32:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

--synthesis_resources = cycloneive_io_obuf 14 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  dacout14_iobuf_out_o1t IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (13 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (13 DOWNTO 0)
	 ); 
 END dacout14_iobuf_out_o1t;

 ARCHITECTURE RTL OF dacout14_iobuf_out_o1t IS

	 SIGNAL  wire_obufa_i	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  oe_w :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 COMPONENT  cycloneive_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		lpm_type	:	STRING := "cycloneive_io_obuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_obufa_o;
	oe_w <= (OTHERS => '1');
	wire_obufa_i <= datain;
	wire_obufa_oe <= oe_w;
	loop0 : FOR i IN 0 TO 13 GENERATE 
	  obufa :  cycloneive_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_obufa_i(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop0;

 END RTL; --dacout14_iobuf_out_o1t
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY dacout14 IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (13 DOWNTO 0)
	);
END dacout14;


ARCHITECTURE RTL OF dacout14 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (13 DOWNTO 0);



	COMPONENT dacout14_iobuf_out_o1t
	PORT (
			datain	: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (13 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(13 DOWNTO 0);

	dacout14_iobuf_out_o1t_component : dacout14_iobuf_out_o1t
	PORT MAP (
		datain => datain,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "14"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: pseudo_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_oe STRING "FALSE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 14 0 INPUT NODEFVAL "datain[13..0]"
-- Retrieval info: USED_PORT: dataout 0 0 14 0 OUTPUT NODEFVAL "dataout[13..0]"
-- Retrieval info: CONNECT: @datain 0 0 14 0 datain 0 0 14 0
-- Retrieval info: CONNECT: dataout 0 0 14 0 @dataout 0 0 14 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL dacout14.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL dacout14.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL dacout14.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL dacout14.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL dacout14_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
