��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�c���-w^�h��T��6�e�z�x�� R�I�����~���]�?;�A�%{�24���-��5��!w��ͧ���x�aДʴI���>*޽$R��Bf
�C|��)G1&mv,)�L��a�\�!�}��h�N6E�j��1
�f�����@�⬼��������=��5b���"�h6��ŔO�����L��0�"�P��&�5�S��-vx��|eܸ�iB�fTV�n��mg�՘�� �΍��� G�v>���h�AD��Z�iڥ�5�/��F���2c��I����m�"�\�aeo�4�s��-�z�x�ՖR�;�5�8�e��?���1��,z�*��N�?��Ⱦ��Y���2�I��=�~��
ɒ���N�"��+3��X��
X�Y���A�Q��I���"0�˼�A�`�j%'j,O0��P��o\w��+���~iS�|��C�������C�^>�S��d=j���%g<�˸�Aװ���������\r���$����/d��%�������@L�}����h'�6��ܟ��K1��.�/���g�QR����l��<�$>��%uVE�1�Tŧi�1�~���l.�y�躪�������_����9�n��i2 #A�<�ȿ���� ����6��G��9���ҧO�0����r��p+Og!6���� |�F�on!孹��XG*"B6-$��Ja�o ��T=3r��f�K����ݻ(�pK�`�����_��c�>>���G�����azR滳(xJ_��lȅTi*0>uhG��� �Р��R�:��*<�i�V���^+�<܏j�?���WJ��u*֥V�"�@�pE�H���������g�G�}BW���w0|E{2pW�n`�%S��˝Ą��]�pa���<������c��K]sQŨ���AT�GP�u��w/
�U�&�������j��9N��n�����0�c7/���SI����������7+�2�N�"�N��Ÿ���i-&���_��}��q�2�Q� 2e<aib�#��}�/��y��6S2́yīyY��I����8 VbK�Y-��;�:C
Ƒ�R�!���T/�I��
x��Z�L�u�A1x�IL���^�!c��su�����O��Pz����k�I��9rl�I��bW�<�/!_��س��n����t�����dq�f��=�؎@�N�v�\` i Wl�C�=h	�b�Y�,�{ P���b�,��|�v���5�ˎo�)M� ����fwS�ש@���'S˞�'�R	w*��[�ͫ�Fޣ�@ܨ�Ǒ>ɓ��M�5���H?]���Uf/�[���H;�#����}��)�H&��~f֑%��qFAue�kV1 ��ZB���8�6�m;l�A�_`q�Zfcx1^y*�+ �/�*뇎h��~�E�Y���d�.5�xh.��@P��c�8)w=s(��no;�ԪB$�FI2�y3��Z�*���6����b�����"K�}�m%�u�_�>iuք�g{��y3�ov)���M[�DT�x��d��$��Ig�}�'�����<�L�Մ��~�4%a�G�܆o�5;y!�UM$�&��g ٱ�E�te���jC�F�|gY�E�� ��`Qt�[J@��G�e|�w�ϳ�CL[���+fK0\�&G�_���R�u��16�@9�>'�o�~z8O������Dծ�<���7��|W�ɱ�Jֶw�$g��ۮ�&�q�H�j��+��w�:QKފ��p�_�]�}q��i�|�ӥym��Z�������n3��OZ�f�n�P":���}��q�}YH̃Fiu��y��W+�  �Ǳ��_�cZj������@"S�Ag��|8	���*n*��8�S��.V���VgHD���v!U��%"Jx�_�o���b{:����s�7SVX��b�0'+��vr5�wI$�l��0�68j�Ȇ)���b�<I`Dbr-|�N��O�׹���Y%�=g�MH�)>G�lՏO���B)ڏ�t�XTջ�N��;�Dw؋6)�!KI����Շ��0-_�e.otǏ&$٥(\͞��I9Ǵ76���܄����t���,�'�"�G�y���5�7-#��L�f9��	I<��q��5��;�������8����+��d"��\�DQt����� �W���P1�c���f��a��"@��2�,���5/N� �+�y[v��� Cq���j��:�BW�f/պS�3>pR��� (�^7�f����c��I]�k��	��pȓ�2_���9�;G�KZ��O��k[�mV���m���vq�B84�����W�T��h��GhfduO�۠X	ߜ,!R%	�p�p�)�I�����;�؝<j���I�4a�Џo'L�U0D��t�R�Gm����n��}/b�K��/2�K����ޔ�r���h#�#S��;�������/k��M$��kb s�y��MK�Id���'<&�{?73���D��w9��J3R˟��.E�8Q��������<0�Oy�)�X��ڞ�`yE�0�&�O��!����:5:\b뷖�����O�'��:{����f�b7Kι�����@�����o[:vˬ>M.;:��V@X�Ѱ�pG'7~� �H}�t݈?�������nOx`rsb��H��sGE�F���}'~��i���Vj���0ɿr{y �G&��}԰5iJl��f�@	�������e괸V��7S������t�)�b��;o���ݏ2!�f��ִ��<gϵ�5�1�@-Lh���;G�W�c77U�a�I��*�׋>>r�҈�-٠�W|�<�RAa_}���JE޹d��bQA[nR� ��e;e���K�0�5���<p��b,h�VT��1����j5���х<���Um�:�Z��X!s({��,a��X��a��,w�5����{�塋r�f��!2W��=%Z��@M��HWǅIn[5�e�n(�t]d����S<+�Ig��֤��(Q��|�lF5
F�<�����V�2�j��fC�mfj��1�Âg�jF�.f��Z^)�ލ����$�4=������n��{��)$H�vH�&e {\G��n߶��;�D��gݢ���������	�X�؇H�2`qod�Gh�����S|�F�؇��F$�� ��u�dJ�с����U��ߘL���r~L��N����	Wؙܾ��4�[3	�<ku��Wф�I_����/kD��ιl{g�t�bsΚ �IH^}p.�b���,�i��v�Mqc8�r%����BO+I�iͅ� X�c�E(�&%4����O��M%5i5��/t�����]%>��x1&���:[7��c�٤�2�7���ҍEHz~9c��$�w��$�0(%�
݂�SO5�|p`�9Ԟ[�hZ*VB6���,*�%�M����|���"4��d�r��|ٻb�`�Ӵ�`N�ir���a@�N���N21�[p���}zi[H��M�&zO�榨�'d�t�'a�k�=���D�A�khX��>᦮�8!��U�B]��*���~-n���J�A�`B�YU��ٻ�餾�ޤ�������n%w� Znm��Z����?f���P^:;��:���,w��*�.����pF��tȆ��lbKnʘ>�S�D�9��l ��-����*���ې�s���}#wi�}�%�NG)���Q<������ph-�GI?z|�����оH?'�^ժOyO$
�A|&a�����Kӽ	����D�����#�r���Q��(wx�&�e�xJ}	������M��统��P��$x9a?��W���޵�V���7А�����Ŋ�?fos/�����t)o��ƣ�,֠-C�m��jԍ��JPm�c�)y��+>�.q�B�kN�ZZ$�\;cI 5;��k�'�{�Ž��aA?`�q��r�`,e5%>qٺ�&e�� �A��R�J�rf�N��(�?+��z)�V�c�ӶZ�������ܛ��^���ÇGE��pw�lU�:�)��;�xј:����nm\'O���h���ȷ ��>Md���t}���{:6�x�i0�$�����ǊiHE�yM�cf G�gw:"鳮O�<�Z����m{i��� ��4�ʲ%���U/�'�u�s9��q�.i꟬S8��f�`@wz_OR�ee�ɽuG��F�<���h���-Qp��%F���{�����CW�n�V��kd�8/�ׅ�r)J��{��`�n䪡Hlc��{iJ,ET��*�����
�	�Itiǋ����d.ӱ��J2l�*�f�����>��������]xi�+�F�f4A�r�"�_w�*@U��{6�c���5oM*�f�ɒ"QloLJ���_1��Y<��Iqah�e��,3aB ���W���+X��I����^�����lxQ��\���3�I��h�]���;7��cP��$e�����r �#QHg�͋�5i�@��u�ϼ4�i�u�����}��B�#+���mu^�g��x{́;Ƣ�0��Ƈ f�;�f�\Z=PlԵ)��~#~+B���:�Ҧ��c�dأG8�z�Ԥ��:��J�ޒ��3�l�D�Ğ!��e�������r_E5kk�户���{al�`�A�3�̕�?g)/�\d^bu��Y2]�QeH�@��6G{1�p:+��B��'�A꽊��$���R�Hy'@��.h��-�9�"���6���w�B�`�
�|��`�|7�%,� �� T'�+��?��MB�S�I{�P7�VYj.��U�[�4
�t��.��ձ�`��	�\q&:/��m��=�(���V��9*@i��v'y�\�s����}%���v�}-&���G���>���[Oc{T>�~�Kٱ��݉:��b�7+��,�C��;��"�faK���z������~�P�&���ޮѰ@�&F�|����xMzR��9��r�.0��� ��b��5Tj�K��=�O�	 ���oƑ��f�ω�Ĭ��T{]��y9�x��Y��͏����P���Z���A���S�0���);�j�\�4xs�}}��
|q0Y�h��(��?���_	��	��*:����PM�r{Ijoo?�{�]/�����?�d�,�k˟�YFH�MɇuO���,GZ��mt�E�	�1�����($���´^��2��l�Lݎ����>׌2�Û�z�o���=( ���V�7>��u�X8�
�����)�L��R9�_]���Mr=t���%��^xä����mdEL4I����
d��riLT�N�ݎ\�w����fa/����"�h��?6�%�FvX���B,<9�/�F���=���� �����z�t��?�?I��W�9ۙ��mʘ����
�#i��?5@[J����B�����hk�Q�9au�ώ	���
�4�L��?%<�q[��@6M_�k��o��14Z�P_�Pd��5ݴ,�@6o�L��&����S�M��Sd��$����w#��
4���b�:�U�aD?(N{��X�O*���h�H��T����~����Ձg)���(ЊS�6��p}�L�_��E����o4[y��9��©��?��r����<�á?I���/��>����Lpը��g���)��u�g��ڝ�bKV]���Ar ���YoŐ?��_ֽ�"�k�A��=g�	2eį'��(x�D��D"������v0k���F���3�`��t\CbE8�pV�W`�QPrU#���<�.J��1�ύH@��߬�Aß̽�D��yc2��b;�i��Z|�nP��$�t�_�t;�ؒᶒr��ţ��J������v���+.A��<9v &�{����b�����E9 	��$9���3��9�%���r-���C2+1�?\Z�l����
��F��%�u�CD�`��%��vNI3��8Ff+PeXVlm�' �2d=���^��4َ�!G��U�W�nf<%���G�;�����ݤك���կ3��^�8�j�"�zǖ)Փ��a)I�x�>1�|sT��{	�6F��Z�F!��6y��4�EJ����7� ƍ>&&		�~��J�������G��Κ����!��+LZ�O�
8��Hn���q{5W���/=:c����^�Q�Z׺�ÅѬn�]E�R ~^�d4�HHS���X0�3��F,�`���M��`�#��ǳY,i�8���ݍ���G:e������ݖ����eR���A���f�S���J��FH�i_s�x�?+"��o՟#a� ��Q�VA�9��?W�BD�F����+.:�5>`�{Q�W���h��	4B��9�����W�OEҘ1�@���\i�Q����x��R��d��Y��R�C<��h+�l/�1oG��	�Jǫ�l\܊.�Ǻd $���Y�f\�Oٗ≇�jݫ�Ǻ�\�� �2D������v��~{���b_O���uyLG��>���v���� �j����`����
̃����(�}�[`�n�\4��S`+25[]���_!DM�S�a�m:�;��tx��*�sG���V.ƚ�.���h�ڄ�rLrTП����m�ҍ���F:.�v�NQ�QC��t���0�͠wDNN���,}g��)у[`h)ǣ#9�\͜�������ɓ|.U�"I4��k�)f\p4 �W!O{�r��cO���t�1�@�+��[�����LL�������,�N(ޅ���C�5������FHI�b��[Ԏd�ƄeIx��1�~�W`�o���s�Y"f�u�����*��-���'[�I�҅��E���R�ܺ�m�r����f=��yh��żD~�&ٲ�;�W��b�<��*Lf�Y[�2
��\���B������ ��7�ҫ���r*P���9Q>B�O(�����x�4,o�& ��������9l�*4a!�ړrNi="�*سP)�o¡O�
�u��ϘׇK�d������O�(r�ΥiwiEv`����R0v6*� �eL5v9x�Қ`���y-)K��h����_�Q����tqY�#���2�4�)��0�ڻ���W��O���/�poj_�H��U�H!D�'\)��;��Q�KO��VY)�yD^�~�o5c9��Ơx���R*���leI(xF��x��"����v�:6�K��W&�&Pz��O�a�0��DM6��FT5�ј���b��'&�3U� k�;/8�qU֑w�C��"�}�tx��*�EٕZWS
�=��'HX3����떠������޹��K-�����k�t����1`X?�Z��s�5s�fem&�� �Qy���B00[أ��K[��t�+i<�Ѡ�	��g9CG���˛bՅ<!¾���#Y-HO�И(���1���$��*^�@Ą�[���J9P���(b1f�v~
Z��X|~�3].x��M$��v�Sh~�y���X)R`��Hd�(%Ұ4�m���/!扇�����V?s���F����u�4UgUܽ���Ԏ.9�c�˛��lj�����{��HX����?+{�N �?7�ĽC�.ԋ�^����Xa�KE*����Ѫ(���j#�ea��~�㍇E(���?.Dx�� �Ys1D�ke�5�Qe)[��۾w^=IN^�,�W2�c��"����fMQ�¾�Fh	����/�	�Pt�՘��^��ys~ҳ1#/8��'�i�XzE�'�s�FؒzT�������y��B�7��ၱۿ*�?s����-�x"8FW���r��[�:b�y�祂]?pW$L�Y�_�&()�Q79�|�����^;VD&�R�ɭ�S��|3Y�}/o�C�J9�� ����빺X�5��CkUK�S5;�C�Z�*�~���R��wKD6a��H�{g������5R���)�{V5��Y������E�)�ɗ�ȼ'�l����0�kw�Q.��/ӛ&KH�+���"�Tf�@:�x����~:�Z�~������
S�Ĥ
Ƙ�82�P�z��ĩEm����Y���>s�;H-�$���*j���t��I SH����3�m��fj��6)�Ͼ����iG=|�/@��_y(�b�vzZ�H�ߐ
����)>�+}a�@ v�ib8%浾v�IdQ��[g�'k��k-�kfX����mJ��Udޙk,��Ik�p39�ǅ=|eם�7�C��j0s4������9�f���X��,9�.ʼS�^�'�}�L��3�����n�@Z�\�vZN�S��m��p`J�e�#��O���c��i�T�fM'z1.;>�#l#��{������7g�%�c���1醺D�mՑ1�>�d>��Y��P�� ��͡́�y#�@��N%
/��4gtf�r���ѹ�*.�o6K�Y:ˣ����B%�
�.�Н.g���*�����|i9��>���!�C����=�˳�u��9H�1�ehm;!��JD���9��Q]�Dg@H��*���6��d �ܾ��lX���.�G��{��Z���5j��
�^^�˺���a�mA�(Zɞ4� ��_d���_BU�t�%�*�X׬��mI톾e�za�`4AJ����[��(���æ����6�.�*��MgrY%��~:���c*�L�����&ey'S _�N�_�-����mC���tJl��GFk=g�Oq3��VBA�D�G�N.>�Ijӭ�eW�X0�Y$����i�\i}Ó8m*�߄�r�k(-��zV7İd�Cg�i}���/�f o�[�pr�z�n���у��b!n�أ߸�	���f�@>xB-���M�`%=��b��oJ�����Q�-dZ�^Wʐx��+K�$̠�4G�q�F00��o�x��E��g�9̨}�ރ~T�pgՏq�yL�T�Š\ƿίx�� _�!��^���R������jJ�?5��Z����	�z*� iD-krK�>�q��,_b�"-rӡ��Up��M�"� B��V'�(�/]�Z4�����F�x2\F\	ܳ��cSciƝ@V�M�q�y�,.�.��
�F9h?y3򖣣 K��A+"L��;)�������)eS��I� 	5�2|�GD;�2�H�W3e#z�M�u��˴xA�V���at�n��I���MOD��q1R��P+�q	��#�p6���r q���wX��0gl���Ӥ�e%I��5K�I�P5A
��:�}|P���aʗ���FOo���T4�@��T�R�C%r��<1��ޭb�$Wj�����N;`f����r7́%��j��@���J���Bl�E&SqL��t��@{pP����>ҔV?M���01�`+)�Sn�J��dM(e�|��Ga�����^���8#���-��O�/g�SF�B��~�����V��U�J�{@U G	�ɾ��i�E:|�n(���9O�ݢ���PEA����lhO+�=�9z��-P?aoݽu쵆-k��XA��>D �Ӿ/�4xU��y�<�BA�R%?nBn��o:׽�X�Zԑ�@w�6�ĉ�W��!w���"�T�E�"�� d���<;�o�T.�N�DI���U��
�J��0>�$�
�[jt� �pe��-O�U���H���.R
l�����]^����/��NJß����-������з�5]��}"�=O�ç����~_J�zH�D���a	�N��A�{������ݰ�>s��'X��9���Sl�+��]�a"1� 'i�dTZIbO}!s���3�nљ�?խJg�Ͱ�_�WN
L��vyu҄�z���T�6!�z�F�Y��s(3.:TIi{���F'	��:;G�`����~y��vuO�G6T��}��A�ǰ����/]��ձN�yJs�*�c�+_��&�����
�8؍�h����a>���ED����D���â��I�Z&Tq�-�y�]��j��|��K��;�|a�d�M�x
�}�i����HE��4��]<�ʝ�0�U�ɸ���%O�_��vI�"�7��P�������U�7���'r�;	�Ŝ>|ߴ��9���B��d5�����_�1Y�H=X�&�n��0�t���%�_Df= u��0$�}A��U����yaΛ8R��u�z��u�
����ո1��l,�a��Bњ�4��Ên��a�	��!��&FeCWI��6��"�PM;�lqH0�u
>bP!2�I���6?�X��;;�$]9�^�~TP	�b�����B�~�XV�����O���D�+{�kx>����,��#�_�����MC|����^�b�-߆\�:��Q�FE���'C�r��𰈿�0^{e4��SM���5㪝�nx[�`�����DHsLJ�eE򞞱�R ð`���`���e.�M�w+�
�Y��>hY�/���04����	�b�X�����[�	�^�^�W����福/�^a|������(S��=FT�� ��]�����pj����n{��M5J	�'�]��4Ǫw��#{���)Ԡ[�>�1����͡��`L�=�k޽�|��bb�L�pnuqY�[Ռ�D�1�iBM��TNl����nQ���E�钼Yk��t��\�h	S�K��ӥ����{��3�N�8_E�۽���-��`3+4���ƺ[!�H����p�
8���{��ik+�-�S��+E�]��'���(\E�����ΰ���dȖ�Ԣ9~Lo�Z4�E��)!�֮��&�2ܺg2Q[�ާh�J�zgo��f~�8����-����R��5��`-���b �)�%��q�Bަok�4o_E�	�����H/�A�I�ݖ�7�ۤ+ʫ$�C�iuRT����c ^>�럖CG�s�AVw�I�8�h����{�/z��a0'~�p� ��=�+�O�� X\.��I�S|/��Ω#^df�Ȇ�:���{�����ghX�nޣ����7��e�'�!��cvx\ľ
�Y1ն�;�P��`n.���Y<�W�s�#I \���e�8�q#.(R�M�}]!�6^`�-��-��uw�:��"��"^����WO�\�Vѭ|+�!�Y�><HQEK@B�����]I�f�� ��c� ��m��i��`~��x�+�I�G�ITQ�5��;u+:�s�H[���A������X ���#X��N�6u�`��:�:r��6��(�9����kh�F8�*�R��L8����g�icR�/����I)8������܀�LʊI�u��a���d	��8���0���"_f���b�7��v�]�=K���ׯ2��Y���1	^]ԕ���ξ�ػ���z��&	�Ř<NIIzP>�Y<AYe���ܨ��{��܎Ux���*�lҐH�Ũ��_��4Ω��Is���"1����\#�o>��r��< .������y��!��߬crd�[Z( �R����Yq�Cx3��\od(�VH%���4��y\w��w��o)��6��bj�mP�y�k�ʒb?�i�я5�JȬ�\W|����cLW����WD��w�kK6{�x$�da�`����Fy~P�%�F���A��\Rj0�v��~~�������em�-�x���[x6LA��roF���
E81���I\i0W��S���@�l^����+_o��˷Cյ��,m��.��h���v��%��)]V���#�ĪѴB�����$�F̜C^\h�BF� y{�D���!�5(�K�>�z�N�*g�x��
|YD}����1t��j�c�a>��E3����`Iwn^�v�ʉ�L �Z�v�xZ��L?z�;�WϞ��:��c���P.�u��I�_E��x�5Gށ�-jfY
��`Ζt;�F�]��CM�Ҡ��׊��&��4g����N����3[?��5;����=�`��Ң�(4��5���3�D�Fȧ�'pƦ�C�*BgR�^��BD(x�� �Ds���t(�����K�}��r�����w��x3��z�C��i"����q�dǉ���������S�"�(@���������E_�ػ?Ylk��Z�R���_���x�6K*� ���'>�a��Cb�r�ω5���✛��Y
�6;�1�����v�k9@UGt�X݊�W��1����_�P;�-O�A���=M����+�jyXm�t9�$��鐀ɳ�Mި�W�1����͡M�%O;�8�����X�}����J�^�#y8yh�U����g������0+l���v-S���.�x�瞹�nx>����Z4��uz�ec��a���q��1|������O��������؝f�z��;W�O�>D��fC��9��;4�,pg�4|W=�M �0�����"C{�B�����)ƷrTi���)ZuvE����-)獡 q��^Џ0C�f��$��c��T9�F������]�tO�R��Rg2q�;d��$�׺5�AWst�	ɻ�
}�$o�w��*��o�������>�4qO�W��.L���u��q/�u����Dh���?sqW�b� �/Q��T�)$��� ����@�`�_Ȍ^9����!�P�_�� ��� s�K�|ķ?r�&�2��m����F��&H"*k.���9k����y�t�|��fw�o�&uY�a���{ƃ�x��ѱ$Y���$�P@PLT	�h�[xNK�+`
�v2.�<��_ L����Ѿ��J�x�7���6O�?B���S)�7����3�<$�Y6�T��fa��I<)yz� $�w3lߕ��:�r�͏&6����muʮP뼴4Bʚ/,<b�'F�?�q��E4���E���8��K�$��l�B;'�QN%駸�(����P|+=����
J�	��L<�J�؎�x��p�q8K�m�ƚ|z�j���S�=r����������N���6��`y�3:�=ʀ�Ch�9t�T���Q�ۜ�[�ŅQAT�'��[*fuU��i5c��~���UIWT���9��s�"ܬ>U����_�j񹧱�ԨjØM��t��è㬳?=����鵱�(��B���Ꮆl��fd��Q�K��
�*����>���Hݛ��K��ԥ�(ӽ�T��+=����fH�����wc��ɥ����8�ܚ�H7�!��_�������Rv�
�� �j�VG
�&��������ç���\O��z s^��S�����v��$��a5. E��� ���Ә�vV2c�YV��=��䅉��sەw�GEmS`3ii��8jVO<J�.���\F8������5�=�bpZ¨`� ��=/t���N��t��?���B8�Q6�A❽ƀ�������$��?Ad�6[o!?8���k������eG�����]��j�M%V����ɱ���=�0�����{��M޶G9J�5����Q<*�9:�W��ږU �+gv랯�#_Z4�nF�*U��L֖H�%/E ga�/�.��$/Y�*fF�yr������K�T�b�����ۀn��g�Ĳ.�Nnɸ�d�Ꮼ��g
fO󀹷�t'&���A��%�ba�e��;:��ZwiZ�f��F��&�H�-�P�Ъ�ɤ� '�Y����,��<^د�ڭ�8�y��-�������Ό�Y�f6���c��"��=��z���~����6�rF\KD#A�GJF�T��ͬ2c�8P	D�*�� �/����ƅT����3��l�{hA7��������I�.�r��W��p�*Os�S%��L ��1���⦥�Uݶ7[[$T��v&�y��am���Kf�l�4�?�j)i�A��J�@�½~�m��W[6O�7�g\
�o��Y�R�F����ڸn��0#�ȳ=B�K�wu�(�bW����O��tt�
�O���b�!��#��X���5{�(!g/�F$���(��Tq7��I�0��D��ơ����i3��G�B���Gl02S��ľxo�N:�mF�txݯ�S����		X��M�76OB�;�{���p��ˤ;���"��K����nE�0f�f��7�Ѱҗ;;��4�|/0���w�ڬ�ˌ�b*����*q"}^q�����騅���j�^W�eJ�� m�Z�^������?{"_=�#@�����GI�����z��F��l�t~[,X��\��b�*��P�D@���o-�XP�֍���=
H�"7�B�%�sb CǊ[���+�;d�y����d�^�h��6�ؓ"Qd�wPH>��J�Qy��"�o�-(�`>��eA�J�t�LPyu�O�~
qQ����&��j�o���]��1~^x��];b�MX?��|�4{�����a4Յzc�Uo�.����1��Ƞ��p21-�Mti���C�v���DU9���A�cN�Y�U<3�mQ������'S���#Xp�N���h̫5��ǕzS�C�A�q�:/�V�<zM�+U���jD�J��^�h�Dr�������ds>&��	!hh��;M�<�;��.�f�w��!�Kw�q�jLc�R>E������%rɇ��S0(7��_�m�!�$%4���GvTZ�X{�Y�<_�����,��rL����$�Oċ8�߂���h���V�ӂɑd:ʣ#�7��czM�p�~���W������)�����/.	:"���{��nt7�:RD�k`� Y�X����9��è��Z?�ΌWd�]��z���+�a[��d 0<3�)$A��h�kA�&���%���Z㨧qZ��(�����W�Y��gМ�h���{�*#I�����$Wąd��Dk�	Y�	����	e<��&)����������v�>"�mw,��d�ttM����W��X��ň���"�ޔ�g��A:g3��58�G�����p�w��YZLiD`@�&�r�,ؿcO�>C��d�]�ʡ�E*k��D�M�;�3�.���_������`1`H��A87���t\l���5�;q#C�8H̎g)���t����T�Z�1Rx�6#�����t�#������{���]Z��ސ�T�a���B���	v4x��Ƈ�WvҀ@#��\�צ�L��BQ�飾36d#-:mPO�<k?0��d����ID��n���/жy:ہT/��rG�vm�0�w+���]A>If�V��К)�*�P��yK^���ʤ"�	m&f����)/�!�8�����|O�pq����*$ė��(�8��l�d��X�;��栋ٻ�<���c�����#:I��am��s1;ho-J\YfB�4��C��C�����H5�A���u�h��~'��z(��5ho�k�Y9g>,^���m�㺮��I�����s�$�+ӊ\��՗��q"��,�][	FI�u_��X���+�����¡�6�5�����D�j)� ���$ �O+�&�\e\u�q!��%��n���&��m�����H���{��A{(��Y�J)��#[�3`��H�h��2M��V}�;�ӗl�
�2�15Q��l,3��1�.ڵ-���u1��H&�U�u�ůP���Iۭa+�3a�qW'��	�� Q�r�� X�Z�=)"��@+[R��c��t\Q�Hk����7SS���H����s�'�չ����4k�ي��׀���d�vOY�j��栧_�l:�Rc`>W	@�ufǹ�c|��((&�@ލ��w��Ȝ� "X��P�_�4ћW63����U��͏���!��o�������kS���'7�W�U@���c'ҿ����e܀��""zh���[0?P��㯚�Ҫl&E�0�4�5�tk9P:;
Re�?��J5~�2EE�J���� X�
�[�p T���k�>�l�1ꓒ%������e�/��mp���wCw����k'Z��$U�Ic]`\�l��m�E� 8j-��(��,�"K�0��U�n�n�}ٝ�����$�>�� sP�S`*3�;�f���Mⵒ�K�ȢWF�s�?�n&Dn�Ñ�E'���s�w�X��k�1���%��8H�������}w<L��/�+Y!�'���O�[��i�\BwL,��۶���7&d�CP��\�no��~�b���G5��|1� хȘ����M�·����¿3Cu�FC���<L�}�e$���H9�*8��ۢ��6,�_���9l��@��S�I��#"q�KeM��4�B��lG��)*z�[[�,�Rv7�&�����@�ڠ�R���D,�d^D�M}���L�,g,,7�.�0�J"o�$V��LP�j�caW�D��$�Z�=�B�ؤ���X����t�G�4&�#Hn�L�T��Ƈ�	�-��ƒ���g5��>D�Ֆ4�4s��c\2�<\�e&�Ӱ�v7������0վ)N��XVV&>�0��H�pw��L�cڊ_��M4�ԭ�g�dN��X><��hEL8?�\܅?| (�h	Y�ͻ:B��eR��H���Y!d#�k4� g��ƋЕ��򠅙�:�[��L�'�y�+�qu�L&��8�D�2��P!��!�:��NI���ȭ\�3���@��]|������m�H��C��[eNYi�s}�S����}>��7w��x��m:p/=A�\:�A���p}�q���u�i�n��~D��~�ȪPM ��t���=.�@+,oH�������]�&�����^U�b8�5S+�
pv��͆i�΀����.Q��C����4�D�@���-2�J�����X�:�w��e��S�b��~C��-�α��mY�8&��=ȋ�K:�nL*��g�6�*�";�k�"|��It��SkO�LiHp�ͨL�zm�c��a�cjN<�w*�3�?C���Պ���V
�ڊ{b9����i�Yr�A�u"�2qV��f.BıԷo6�a�7��Ȱ���S���<�a�S?��5jxR
7?WD	m!��)]9�~���С�Yؾ@
 �c�G�6��5,��Mj��ݓT��<<Y�øK>���5q?����J�<�3�`���,64�'�v�z�!�ϳ���l<�.����$a�0 &�q"W'0Fi�����-h(�@�� ���%Fq ��F5
����톢�s&Ee
���d�_�6����Y�%I��Yx��og��A�\_Xm��c۷�49�{sO<����P:o���%�S�9�S���rXƸ�PSv)g벓s0�rEλsBO�~뵟P�c�DT���|�D�50C�Ӥ%`L ��]*�������(�����6x��h��[��t�L
����a�w���c]��q���Ƹ���襾h��������v��y'�c�9u�ԏ�u����,�=}�ڱAB�!L�N�T�(|���b���0����N3fO����q�>4"I���,Х�L�����5x1��̳�Jm��1R����{s�g�~3��
�����T"�y	(���"���>�"�K��k� Dِ)@@�{�[�-׭��2ԲV�JkTB�h���%���IF������e�D��A��
gҖ�3��czڮ`�����Ѝ���o�^����}����&�4驕�%�	��0�V=j����>MǊ�w������@PC�T���}��*X�T_�P�j��2��&�8Hl"�k��o��t��U�E�����E
c3i0Y�c� �Q>�PU��;}L��Ћ����?�דH��|o<�(;�	�����ʮ��{hN���Cb�zeU*��.�C�B�Nʌ�Q��ld��Ÿ�:.�<�Rco��ξ�Z���==���Eߌ*��Emc{5-f2���״'�j�ԣ��Y�2!4��s^�C�k�ʹ��X�ͫ�9�ɒG�OX}R�#[�:��&|�t��2�!�t8_�u��6�T-Θ�w����������`�ܱ������)�U�j��2���+~t:e��b���|$#V>��2|=ui�7��D�F��&�|�fJ.�T_�i��H��&�_���U���&��U��ϼK���uof!#���\��wс�Tl���ڽ���x�M�����H�y�{����Wa*��]Cf��?����d�<$���n��!k��q=�j�Q�P��C���;�IhH�5��J�&[+�����qbK�&�׈r�ޜB�^?7x����LG��J-.���'�:]�1qFwi���l��Fc�$}#��k�A%],����`���V���G�%�d��!�W������ �iد
�^n�ԨZUV�Y}�e��74�4}Ս������Ktu�9xs9ρ��8"�v�`�R]o�٫a+�� H���п��*�+��]�aH�C���[��2n��q����Zx��!�֝�3_�WV����o�������"@5��ǋI�Zh7��� ���K�z�1��S%b�nk�28]�K���pa �sҐH�8�3w�M�����
��+�xd-�j/�=�
%�}�S$3W���&����)�0
�4��@N@8���g����-�S7oJ�C-��#i��ng�4��7O.}�?hij�H�Nۡ(9��ϋ��FzHԪ�H'��>�V�c�!�D�lX�[���0ޣ}y�`t��YO�[��r}vA���x����p��&ħyn�	0p����p��a'k@A��tHG+�/��t��.<��t��eH�qY�F$���Z�����$7H� ��o�<p�x�~��������7''�3� ֬$0$�D�]y)�����s�R����:��ȳga��A���؊��M�Sk��2� ���z��+��ܜ���zv>^���aw�yN��xu_Ŕ��~k	fK��$�@ܸ)-��.<-�#\]ru��nB�ծ8�D�u��Fy:�3�{8~����.��3#��)]x7���7��x�6"�L q��3��l�2w�o��L��#ލ���T�K\/�K���~-1�>�N{d��M`�b1�!=>΀���&�!���Jm,@�����oz�Аz����ON�5�k6��sx�IW�+�
�k���Y�՜�q�x�f-�Om*��5�eR�$�C����YW-S|��qѨ�_�d-v�X�L!�DOf��(�'��0ބ�$�b�%V����FQ_ɿn����ܝJ��uoO����B����]˸�벍;��ӼR��V���)�wō���YqU��^�Vk#����;"�M�#��M��dׁ�w���@Eu�䀨 T��:��.�a{�4�]QsĔu�jsp�����#"�)�b���ܩ&�(ԸmGu�=h݃�VJ�S�F� ��֛�e�����.�|�̷��i���Q��@>
�_[�T�g���e݃��\��O�GP �Z���ppA�g*��l�i��ò��� �Z_8y�8j�]���$3>���7:��z#{OF@Q��!T�GKܗh���~�0�2`Go�(�R}�U��h�R_���� ���{	�-���L�P�O%{:�mr��<�ݘ.���v�7��6�&�V�S�RJZi#>��g3�TX�#���.m.E<P�F��������Ń���tG�7G�6Wh�r_��̲S?���̾�*k����0��tם��h?�P=s%*�!��MF����m���PO�.�y���Nv,v���>�5��>LĒ�%EA槞�4��$��2��
4;j�(��o���0�-6A�F��p�Bp�w���O�7l��e��<5CIA���v!��r��'dN�4��_�����~����0v�5��������pM����}{/Y� @B熸�7��3�LC����8������Kx�Ҳr�s �t=; .)`���sS�;����k�1G���/�:M�Ǉ;���7�~��urO���~7���^��|��Iv?�2�=<nd9�#��`����)[a0%���>����4�Vč����s�8
�qv#i{�N���!�[�����+�����s�'�T�76W�Kp	S��Z��i8�y��"��B�~5�Y�7����<�	z�8��lSG=��ev�H@b���>E�`GdW�.G,��5_��K�uޚC�q=?�9d|�)��L�E�`��O���0�y[�Ո`;���zs�WWE|� ]J�9�3Ѧ�o�tO��V��_��BL�@�0���HK%����^�#��׀0�����l)��&^?*�~7S�	pP�����h���'2�cU�wyi�B���I�9�����Sl4i"6��V5��cU1����o�T������O��o��I���I^�~,����h��A�-�II��A������9ݻ�V���y(�� ?��í�n���	}�KWȰ��t�q�^�u����׃@�%��R� ��Xr
'����w��g
/�I�n!a�8 �T��7d�(�ڦ�.yK�q��ŕzڛ�k��ߠ��6�D��=?D��.O}�[=6�&$vv�:u��e�R���7�kvd&�Dv�<`P�_�0�GU���Apᘃ��U�Ŏ�/4��ھ��J��P-��2�4�f����������iqM��Ċ�0R��1�ZJ��96G��\L&���K��'���U�����;��j	Մ�W�i�AW��8408�
z@E��ے&���.�M�f��&=�a܉r�Qgι0��5QX�3�{7H�a�Jx��2���F�������u�|�6
��Jw� ��T�秫�3�
o��������N�:�Lr�_��JeE�i\ь��U��.kX	��vi�k��b^.�(��$l
�W�N��L-G��䥾�6���1�����Ij'(z�Kwh�q�{���g��F��I��ֶC�.X�$�%歺,�vcof���a~�/\�J���\w�p�O
a�eY~�����A��q�k���bۣ�^�h�ܢ�L��-+��h��� V�c�����vz.n�"�mSXV�v�q�0�qeԊ��و�'���@}@y��ak�`XA�Ë1
�,5�Ň����v8@+�F��[������fzX=��zm{���<��S@���r8�G�T8t�7�%{4j/Z���\�F�ݕ��KTx�q�sҳ5��+Ȟ�3��_�!i����ffelbƹO~���{i�G�}����~f��ҵ���ݺ�����Z3C�E�6/�ѿ�-�H�.!���k.�xq�K˩V���� ��4/>��Nl��W�\� ���$O�GoR�6ہvY�Q��6'oP�O'�w:t����FQ�<{�9���J�L&Vm��$��Eo#86~�a���!�����?]��!x>���A�����X�Ӱ�e��U�mp�{�K�c��c튱�kj0��*8eӽIN� �����^�v��o�.��8Θu������~�D�os���A��w�g��Dֲ��D�M��Yx<7�N�>���a���y�}���w��X���Ҏ`j���g�8���[19���om���Z��A��"sƔ@�T�TK�O�ƫ^�X�d�(8���f|8���Ґ�D��\�d� ��V ����4~?�$ ���Zm4��}�S�0*;�*wkf+��д4q)4��}v��\sL�J�Rz��K�t�u^���������_�N���;���#ѭK�lY���^ft|#��m"� ,���n�ǯF�b�Fg���m+�G��s���o���`�uӑ�u�?�4��� Б�g���燾8�j�;d�0���-F��Ԍ_>�4Y��f��G�⩀���(�x�!�(�ryC����!��;�ީ�}�]P�Y!+v�Ĳ�l�}<ˠt¯y��l����=�@}6j�����@y@Ę������K��^�h���~K�<y�Ǣe�X��������� ����������F���-H���!0n~�$�#�(
7q����qaf�� ��5���B�r!<O&��%eQ���78�;��,a�g���ʹ[���`�Rx�PT�,�������x�����Okef"�{B��k^ ?����PE��ig����}$��u�2���?x��?w8h&P�a��$���D�w�S�����S� �p(��`%	M��D�2?���$g�f�4�U�	>'��q��ɼ^������Dm�(�lצ���K0� l��AF�-V���Gȧ��@V=P6�|�P�Q3���1���d�Ѫ�����@m'���v_�P��*���x�׷�9�o6�&G�k*�=�Pr���ҥ�D�5����X������\� *-�S�)��ېs���6:�+��\Mh��vH�7���a$�j5�;�Y*�Zz؂r'B��0?��{�G�X/%_�1���Q_�%�Q�'X�FY0�"� 6�N"964�*�>*1$���\�m�a�� {s�y���L��\C�8�Jv�q/݄=��f�}�I-�oy��"�!�N^"�n$�:�R.w�@���g��;8�^�T�M浤5�/���Ms�|����5����&��y�Ԣ;�j4Ch��_��Zc\��9e|�:���)�ޮ,���� �a��z �	Ś#�����kD�;�Bp�Ċ��!\�:@H�Q���3�T�Y��*�.@��ѭ����ro^����$�*V������$�A՗�jF�Dq��B4`X;j8k�:s4���:Y^H6�,���)�y����Y�V���r#Fi�'?��6t��o�E�š��ـ�l��y ����)�7�mj����� {�,�����ܕtyPY��Ud�����i����)�r�].	>�v:(��?Hy�C�?A=�N8�$@�|��~ڣ|Z��
��~�qE9[ L9"��-ک�Τ`D`R��\2&���X�+k����M�>A;��+5m�9�FX^�1�ݻ�{��u{Q-Sf!֝��x@)��W��Hh�_��Y&=�Z�K�@2�����u�5n9\�!A��	SR��������N��9���~�:5[N�!�^#aS�Q"��Q\�X�ѧ����Agw�V=�]?p�	�g��(�3�=*yP��@�6��`��+m��^sW����އ�(L�E ��p�<gM��F�1M��иZj��Tǌ $i1�)]Ӣ����M2�g��U��a~
x
 ��l=�̾��p���A;|���_}ru�I���c��!��/�YY�˛wt�^�N=��l���|�UO �*h�-�ѷ2�!���gt�)���D�.�G(`a��/���t�Ihn��{5Vlz7xLK�0��:���5#O�m^	'��VBV�����)PQ��p��T4�F!����9`5"����� �'Okd¢��9L�Q��%��=�_���d\�L`�٩�ҕ��nN��<�M�lq��K��h�����������}/���4y&x5Z\��n�el쌩Pl_�F������[[��;"{�AR�!4@��!����ܠ��n8����ϙ$�H��C�~�P$�1=��w��n(L�+����K5��r��>uG")z�y�v.���]����ҋ�����T42�w�6�ꩋ�DE���n5�z�
�Yy��|��������[8�ɹ0b���_$ߪw�Ǯ��hH���K{ �C���4�+c"�$�����F�ޣ���5'~�uc�t�]U���?^���t}a�Us7D��8~RF\�	�����rn��SKG3q�4Q`��U�H	��\kbȒP1r��2̄��"pf�fY�����a1�S��(3MRF�8� UsҩCW#N c��)���'E�H,�8�
.�go{a�ڸ������o�@G6?�D��`�*<�Cj�0�