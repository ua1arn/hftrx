��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b�8N�b��QQ6��4j�)�E�E.��o��.����
-m�w�����'Y|զ������ޢ�`�W2�)?���	*�o�VқȂ�%#�&�����5�{�<Kfh��`0��(�r(�0=uVܒt~��Q� �<%��d��)��GN��zH\x�q�E�[��-�z��5�~��س��Z(L�S��X�49����ZSN��6�H#Y�e�q�q�Ly��w�+´6����P�K�Ty��~殕)�}5�� ��ӥA�I�J������ϼy��i��Ŧ�Ou�] �(�=J���f��� ������pF�R@^s�������UrJ�1��V���*tUФOo��0�l�nJ^q%$Ï��͍!�f�ߦ(�
b6����R�3�|:�2E��'q��<9K�b'����:H:���v�W�%ry�q��%>�0R+!w�_�C�e(Ĺa�DbnZ�P��D�"?���X�[)Qtq���4��ȟ���!�r��D�L�'H�	��9��C��,P;߂ vac/u&�Q/}k�l �:���/.�?���>�{Zз��{b�>��&0��=����6�h��B|8��-��:ݲ�ϧ��ۊv��������_���ZZ6_y)]���ė�2�ɴ:��d1��|JQTf��5+5}�)q�D[�y��J�Ķ7�T�����nک����^}	����שP�����d��]X=��%�^�>Y���_�(�Ő���{��(���f%4�j��d;�۲'��Z�O��Q�=ɥ�J'R�S��.V,w����S�� �9�ٚ�Lz���+=R׎�6"�%G_Z	XL9�`���/���"�?f��bۓ�(*!��p(l7�����*���!���Î��o��]�
E�~�a�xٝ�Ն`��7&̙5g���%2�PQ��NjE�;���/�0�[g�F�[4+�%]�I=$dLr��xc�'^�ʂ;ץ����4"��,�n����d��יهI���-Zn4��[`�ރ�1Ͷ�+\��^�p�xN�L�I�l�ר�ڻ>���~z[nZF7��]m%;e-u����PH,�>�HJ��0~R*���%3f���p��0�\��Rb���ח2�U�MAF��f,���Ԅ����������ƨ��Vԙ��M�*f�������4���{�����i�'���	s��A�X+� QJp" ��Ń:k	F�2el� �:�ʥ��:�5/r]���Z��Ǔ�m��Tl����o`�5��9�*��%>�Q�?�nk{��_��`"�6=��H�������J]��|������ێ�F�W��o��A�/�1?�6}�ȿ��Zʧ.���bΈ�9K|��_��"e*߽���7������9)i4i5��5��6�*��x�b��v���D�{��C�:;�.�tz���UzsQ��B�� �#&:ۗ>�#h���˼�)| IL{ת�cp��GHVQ�[O�i�W�y*�1��.��ؖ�r��|/���2�݊����vҝ(�T?��gڀ��t[�:�4�[���`��1��4��u�����6�6Q�ꤾ%��X���)L�\&]0�jYkx�_b����4W
����o�?6rH"���4ݜ������<6/��[0����~�.(��^,I7�T���y�t;�]�*�<vجH� �~���+�O
�Ķ�Ӥ���s���\�L[���"Ds���6H��ȸ݈�w�0�\K�D[H���*��=���䠪��݇a�2�?�$,�0�_��Qoxn�8�@�iy�r��d̜4R�����硐�BNVVd��g�@5��BV+|���b��(l���3��<����T�@����l(Yg�clۧey*�\bw6���n4��eË���ԧ�0!�a0�:�� P���0qu���׬Oz���cp���<������"�+MH4@J:�&C��6Q^L�JZ&�N]\W�����<��#8S|�%4ƹ�*��gտ��-���4���2�`o���sf4��"H�!
J��_���d�����\�a
)������_�A�̋1s��$7࿺���W{�ʍ��E4Mb��l����b��K\����W� �*�7�s̟� mH�?q��w�5��d�邌ʟ`�#�_:��`�a��4pm��$  VC4�4A,eS}p.>ˤ6�{�6�4��=~yF�	_Q�a�]�����=^MA�4g�������B�Hf���.	I��	V�R�*W���3�U�eO�=��[����Ψ���~�-�7ٙ��Q�Q���s���7��lM�L@���H�Q���'2=Rf,��xx���ܓ��7��i O:��Vq�&���w�c�}�&�=�8�t�
��Q#uf���`�2C�5�?�wm��	lo)���l ��JC}l��a�9�k�k����C��TB�H����a��i ���)���9#m��+�@ș�Q	��C*�R� ^�)�t0��ڴf/'���J3��=�l���ɔ�����pǯ�����%
�x�ŉGu�rXNȤ�y��=��^lt,&p����\ �e�c���<OA`������c��IF�l�Y��YPn~�8�q5���_��t��p\���������r�nQPl�cK���7�;�}h���.b F����{�RqE��}s6[V�Z�Yŷstj������e���S*����r=\��	s��vg�lϩ�x����� �:r�h����&��&0�[0�3��Q��\����:8��=���^��m�� �܂�Ot�UB�x#9c~�&JC����D=��E��y�ߛ�k2x��E9A�M�b�~�E��gq�?ݗ�w�&���k[Z��.*-m�NOw{�L!��0��r}ͪi/�xj;�+����՘3�#���)dܔ�-Wɦ�D.�_����9mK��"[�<9}�Ό�2�;,�+���s��-�lZ+���Vi�m�p��	��}��c�q.D���Ǟ<�P��G��C�,�,FXy\Q� %9g~�(���^(����U2�JT����c�|�V5�HƯA]<����Ŏ)�s����]O�8Ar�4�-�i��#�1%��o�&�2�Q<Q�������˅{���I�5�)�uo��P�����!\e�//Q�,�F����h��'���/�Z�.���޼}w?�&m$�eM�[�v��1fp��h��`�/��c��jn{{�b��/�T�]���v��ӆ��vK�:ǂk|)�8�XD���J��Cz"m��J�d��|.V�2��B�Oτ����rfOR%6`a>�*_/iU�!�K'�l�����^�pT>��S%�c]�']Do���Ai~��l}�k�#�:x�RŹf�Fhw")R�UQ	�z+�Uj)W��Ϙ�6ꉻ-Qh��W��B�c����5�����j�1�v��t?����ր�����=ߺ�Q��VT����[ D�bu��{���A�Y�{��}^����rZi�rJr ������2k�ʡ������^�]�2������_�6+л��Z~1�M��E E�R���'���q�a��t�5d?r����"�ɹ�~9	�~�P�ƫ���W�d�,l�l)�S2��I���4:FO��]����6QZ�*y�D:�V��nZ�vhhL���}<t������y��kc����T�R2���SZq�Op'�r�sO�N���
��r�L��s>Z�9d�C��U+E#i2u*�v�W���3c��0�bfr�M�g5�i����Y�0̼:�1w��n�Q�{����bm=��No2�C����e>�Z�S�Ԧ咄��Y��tK�JV�g���e����dn�
w2�f�yu9G��}�ǩ}�+�;���=-��;᜸i�r�A�o4���M�b���,�P�q�M��V���Dx�R�a�zk�����q�kV5Q%Z'(�&H�����+�x(�����eN�u
�d���cPfa�b�\�O��2�![,̙���H%�[e��3w��Y!�M��(
����H��u�O�7p��4�*z�y�������p�P��� 2:vqZyL~^Gʕ��@�ʜ����l�����n?�S�T����j#�1���x��-��%�x�����H����>�"�W�`��;B�,�� e���T1?}4�:!�.��3b�ȁD㇉�i+q�1-#G��9�%r��j�d`��#Tߪ�Ac�����~?u��
c��0�Vz�nor_]f�Ҵ唵�ǈR[|��&k|�c����ek�xi.u�R:��O؟��$,)�Nr�R�F�����e�3.i�OyX�gLe�wZ�\P�|ed�&T�`��AuO{���ɳ��,A�	O;c\GlA}����s�0���}ـ���Z��A����y�ݨ%4���se���i���Y"�����H���\g�����JI"�}X���Й�_�nd�����b�w!l�: j��C!��0���_N��+�h�>�U!�Ā��^`�zE�<r������U�B�I-)�-/^�0g8`Tn	5���e�n�Cы�@��.�M2�����l������>�#�07A@9��ŕ��!ݚ��|��\E[t2W����ˮgۗ�����׎��������Y�%�͸�^Q�{�b�ٗ�D�p	EIpX���~i�)�&B�6^�WL]�n�	Ӹ�S3�_챖
�U�7"0j5�;�
:�Ԯ��j��3)���sZYy�U�I��̫	Q�WG�ڂ�lL�t�u�����I����f�2@a��r��y=|��[85�"@����|�9Iŏ	~ �j^XGX"3��{�ݺ��47����CNhI_��!P������KK����?�O�hSن�F]u+f�!EVI _(��?�l �'��ч��!�jP�b�TTt�^��8[#9x�iuO(.�K ��;×{�&�x���2p��~�NBufQK�NO�=QH���A�[5E��-l=��&�&�)-?v�D��M�����������X|�c�,�H��x.����I!����������#���(I-u�J�Ƃ�B̈́0"�(D�z��\V�b_�3P�7����I�N��2e6Þ��in��|of: ���&����Q�(�"��nٽ�J��N|��R�Z�V,2�����j���x����,ny��'��)bp��1y���؛D��6���J�sh�`K�ͨn��h�E�t������
7��L[�2/T��
ʁ�ן�kK��u}��t�pd��t��)�`I�}�Z]�H�;��h�<�+cJ�����-��<SqD]��b�{����䶚^�V�&|�?B��w�,��C���״�I�%�������!�A�ʋH$��B6�TG��в�����3LD���L5������0v2�#HA3O}:��BӺwr�<�������a:���$� l�����l�Ul�gWp1���鸈�%��X�m�.��@n6�]!J����+u�׹�x�i-7y����{��{� e��$אp{��is�L�q���猾V����_�H)��B�l�,R8 ��Z����k�s7u��0x�]�S9/a��%����'5;��&yc�l��8�¡Itr�ᯜƺ�h�2�^��!_�q�6x!�@�� jq�C��%�<�k�KZ���FF�
�X�/<�D �)M�Z@�oK���A��oF�y��>Lߥ��E"�Ц�`K� �,�G�m`�:��/�%�Ip)m�S���]\��˹�qDC�Z��`�/�z}R�m*�.�h�挢� (e���b	H�@�>�Zi�?��7��Ƙ�+q��2�9ni��A�-���m���om.#����&�Y�u+a�8��k�KD�dhY2�?8c��I��>M��5�d�P��Hw�S�g�*�Bj9�ٰ�5��^�#���?e�K��A|��MOM>���U,g*��D�&�˞2�g(��
Ț�1��{tC����3��s�#��DB���S���!��[mX&���X{,.��2dt�O����bOe���O����x��{>���4�Y���BΫߠ�RbIzY_p���0ѧ4��w�����o-�IY�L�t�D����t���$(�b�	�vF�"݃���3K�W���7�Ν�Q��lGjK�4gp�981���=�oJS����V�U�mRjq��w��K��R��kj�Y9��@���#�߱"V�.�;GP���PmN
�A���-
^��<�1��FvA��!&��ѥ:ԛ׺����-�i܊���y~;QS���CA�eHP�M�����譡�/�]�]֙g�̒j�Kȷ��,��:�r���Yg��w���7T��$;��)K-P'�x�q��6�6�7���n�C!�����:�[�N�!�Y��������.�b��sVL�R[�!j���1��E�,�� �3�d(;X����`-�td/�@+�g&�=�E�����
�Y FCy3q�]E`�������	�ꯘld3f�s�Fw�#����H{t{z��u�A�ÑoO�lV�_�D�� ',��LV�ύ����P]���d�DL��,���*�r*���	{�*hV<����Sxv��I�Z��x}�����΄��aR��1�Vu�T�vW����$�?�D���
	���ί]6UL�`d�k���|�)shc=_`�#Y��翨����؊µMdH7@�c��`��}��'r��&����:X�V��k�+Гu\R)C~o���4`6��L��u�n�̺�N����׀�k+�a6�bш�.2�q�I_�CЯ9��_i
���q�z;�&+���eXN��1l������ 5�خ��Ћl�|��48��O�F�ƷU��)Gx�9�Q=����/�y�&���/eC�lq�E� ��ϬjNk}�҇K�+$:��⑤�
3'��6�>�ImS4����鎫^۔?#/ۅ���!��h���3t2z�P��2��Z'���_����-�uID����!tp�=[��
�̈́���k�|o�D�P�39"��9�c/�*(N�DBa,>�73� ��0�e�!3W���f�ؒ�b�+���ܲ���/�p����g�e=��|sGb�q�{N	�|��-�+��Ȧf��G����e�ӆ,(R����T��0� �����+��^�{�a��}��%����毎�K�薝�?_��/i�`ʍa�VUa�$��X^�0��O@+v`���S�(v��m�B;ffYdD�1�j�u8�|3�u�q����HyW�o(��@�xِ���6�7���-�M�J7?o�Rc�����囥�e�����J
�������Q�fE��1�iG������c��O���C��f�(��j����E
S5��V����O[+ۤr~�py�e"�򨧆Vٞ�4׿0X����V�ʩK; �!i_��GPl�<A�Uw���N��Jq�O���.�L��c��dV�H>�\�.ȋV�0r~�?i��*���;D����cH]B�w.���4��fܰGS��P�[�l���U�55Qz*�j({��'�o��b>&���
�'<^L`F�]X���mh���7U�����/��^"����� ���ܠU���������^&dk+��elyk��"J�1>�!M½�H�������Fk1M���U����]� Bxw5�y�q����T�*�"K�c7�t�����?�ڥx�X�\�W<�ZUS&�|��AB5V=B�J�%�i\y���x)�6M�C��b+S�b�W,���pQ�1>��^�2��βxE��x��?i��A�(����_�t���1��&wu����|Tءid������j��>��/�Q$92��v�Q+)L�j�@Z"���9v8�A�rQ���y�������!��	S�{u?����h�1:1�4��^z��EĤ�X�2^d�3�_0�DE�ކmi�x��Ox��`x��X�w��b��<�];Y=#�m
@4��A鬊�#��M:�'U�4��B}~I/�9$}��� �IO�Sf+JC���|ݎsC�R���5J2�6K�
p��F��T��]A-.�Z]��|�~Xu$�.�Զ6Đ���]��K ���k@)��x@�M�s��hh���l���,�c(�)�tde�+'�����A^�\-(]v=�[��卷L����Q;�#c.Ґ�5��G��X+٧r\�Q�E���DĐ�뺣��\�ѧ��Z��4 �j��!�gAl	�CG�Vl
��~��oփ����Ս" ݨ��m�ZD�!s�Z��!�VV��L��I����Y�D��0�Y|��E��w������B���Ә?�Z|���}����d���6|��aA�z�Ao��Xq�^`��Z�MO)L�=d�}��A��g���l�ӈ؃�a�Yf|%���M�S��,�H�!�
��$�pc��x����%$}w=?�l�?�7E�}R��ث����1Z��S�ջys���d���7�q8-c�-;�A�m��O�8� ֶ&}������	��XG;+����/�ʏ��z����@�y���� ��:ıG^:���:��~�I��z�H�az�W,��,�瀁6�STc���'��ꁘ��Z|P��R�b��Q-��P�qr�Z�f�W�E�8Mk��m��dt�����"�0�Y�LŦD��.u�p�.c;a�M"=������XU=Z�/b��'~�=j�w���.U�~8 �	����`��]f�dq9(������w�{�h>���發I�ӵ��f�7sV����	���d�uP�ϿI���+(|�'-/nPx�ZP��g����@ͽ����by'������I�0gx��e�-H������w��U�p{D�q�걻�ڍX0��O�7A���\!�b|��4��N��É��M	y�i�fخ�j��l��Er�H�]�*.�.�_�=-���ti��߲J����d�(��OX�̉��-��`p]:�1�R{Ʒ�ȩy�� %Y�� yZ� ��F�|�3��b��z�X8=�5fK"JJSo(p�2���K�p�hm*��pf-�h~�w��U�����Q[�q�Gl����%�JYnR@w��Q�6��	�r�ɳ�p�7��o��zL3�aN�A[i�`G�P5�����w+P]7����&�:�x!�f�,	k�8�u<.@o�Bq)9}���>�+�����C�� �Q'٣�Ъ�P��e�^j$g�$7�nr�o��w&1o�g\.5�缀��w�<Q�Fzy�(p2"]Ȭ�f�JJ�*X����,)�H�x0��&�  3���7��dS�0�m����=�"@���?�����͘Z.%��0^a��"X��Eyh:��qz�:�⍅��#���Z|��!��\S=4�������rE�ho��[î����	s�%vRh"�eNv�P�����dz�&�Hh4SA��y]Џ�����W1VB�)���M:���4�#U"/�D,?�S�l+UAe�M� ����*��ˉIl���!�A�,��h��_y)�Q
<��v��e��>-ױ��6e����@JQk��r����if�'^�nv�W��u2�(yV���5EŊ2e#q�P��V�u�_�Om�d�/*:�Z� ��ͪ�����>�Imد����<) �a= 7�g�`.`�����0�є9���TW�ND 'P�g���U!��-����R����u���(1�-�Y�FЖ�.���H'�O��h/d�3�N�Ѩ|�*��|�\Tp _�?cl1BO���������͛"�^<�fX1�՗���tzy�`R�B)?�:�����)����B�{?��\ɐ�4/�%Y0��H�g_�#�+�G�g�������S���+��I�d^�Q��1����t�5c���<W:����T<��̬�hen��?{����˼^�lO�������XP�P�x;��(#����`�5��./_�|V�c�"�!A�������\eO���FF_��qk~���o�h�-�7Б������2^^M�%��M�vƘ/Y�ً��jn�:����&�����PK��ڪ�^CQ��طc^R�4��Q�@�B6�r `�1q�����8O���<�w�[��PK� ��	Q���x�|�<�S٠h����,���u^�-� �-��¬��7����P۰9��`�D�T8o|�i�yh�m1.�����'�S�,_�%��G#�0S�/��qL*��-9�ƻ�	��OJߋ*4�2�J �E3��]�i���b!cP�Xղr�	��
�_º� MF���:���d�3��&u?+2��
����S��5����?~�Jp��4R���q�Q>ʺ���Y�֢ǦZ�w��|0�t�c��]�m1FX�>��',�+�ϖ������`ڐ�Ϸ�/�z����H�\����D���8�u�:ꯣ���נ'k�4	�������c���%<��H���#�5��Xu��(䪌�Sz��\Z�D}��0ߡC��F�挴�[�J{s��!GL㳑	�����ݮ�W�La;���
��jJ��1��k�yy��6< �Lk$��Y�ʠ�/��	� Q�肪�П��NY�'C�x�l���4
��-�0��Ň4�i	��D)꧿Slh\h|RV�5�OH}/��<M�<q�Ӌ�����(�A���}�8pեf)�P9����s�N�g��/e��әy���s�&ާu��&W��B���[a��C�M[o�a�R4��[_�$�!E1�7/�l�a��%Gŗ����=A,	����W]TOH��ed'�ϡR_y&�c�l2���� {C�]A�?r9B�3i��PoбH� g��P����@������m�9 W�f��]�m���Za3�=�5�G�]?Hĝ�-z�b���9n�|���&�\�d�2y����d�:���C3Smi����X��m�4�F�1�m5>�xy�Ӌ�1��a���[�U�RCG�eZEH����]��gX�t��U��21Ќ��/W �Y��y�� ��{�qlձ�j��-u���Tv9v�HZ:��m0�,�7�B����V8'�5�cЫ؄�ǅ���e�ǱM�2��^�g�:���w#�Mp��֦��F�pji�894��y��~���0���Ӽ�s�����	�y1=eϹ5�۞"
,�����T�gz�e��w<~�},��Y�x^O�TW�x�>XV�x�M!-��y���V��o��i�2^7gbӃ�����B�`�6�Њ%�M�H��cN�W�kwf�u$���H/Bo~?8$'q7�����I<�4)���f������$����
\C�����T�1*u��[�ny7TYG0yk��)M��t�Q�҅J����\G&�	��$�Naה�)��Q���^Z�6*�!)�9E�'e 4��H� �>�QI�B���*�Wx�+�]"�L�g��<����A��jS��C~	,|�	�*]��g��ap`S�i�}"k���i����+@y@��:�Z/�� T�5S~��o���j�DŮ��n{�]����E��f�bK�WJ*$�3����|2�d�)u=��A��%���ߓ�W �N�N��7U�J���ckΎ��F��fR�������!��\�������ɱ���B�^J/j���u/��+�C��Xv�B�d��V�����)�V��������6���6+�c�Q_��Ӡi���+����=�u�龅tm�t��^ҵp�
����c�=Z�E�D�5L&eW��]j؋������)�T�{Gp`�0 ��2�R�'��vY\��%��3����e�Ӱ�o�{~�O�� ���!Zf: �k��oB�؞�"!w�8�(z��M�p7���>�Ě��/��qO�*�җ�g1��W�ǧ=������0�hv�0!�4	���$5�?	�?��͜�q�_H,�
���j����{p�q�&����ѷ�|�q��%���։���ؤΦ����$�'K�Fw	L7��"S�)n������<�Fr;/��}�w�Ꮂ�6K��6�����>L�V=�9A
��2\�m+bNDe�Pd�eP�1�y[��r�xoNԆIg\��\����'�D��
$���	l�d��ʖ�ĥ�SL�H�J}.�ͫ(���z1(J���	��"/�����j�i�W�Z�{)Kn����MOXБRx3U�Ę+곲�C�W���H�n=l���m�XK�]C7����3&�C~��P��$��^!�X�l2,�U�������h�����I__I�L<�70�(�ѫ�����}�e;�q)(t�i��b��p�kmw�"49p���W�����?��";	-߫+[�:�F�?�9�Ac`���&�-P|%����o��t`�(��M�Rbp�F5�Z�g��j�2I8a�������>w���(���E�ʔ�!�A}ԛAq��X��SE��1Ł��n��
�>og��r7bÒDv��LsX�+�o��\� >=������)�&K<�bd��@	;�t,��9>R��H=��ޤ˄ɤ�wɟE0��y$:���6ߛ��80+�Z��8m̡���<�郤Q��Q���z,�� }i�X�lw}�$��ӊ+4F1�q�f����m�|�#E�q��i����L��T���0 �5V{��F�J�7޸1KÍ��p�1��е/?M�N�k~Uf`��M�����bn�-���s�b�h��^�|hlL�С�Q	�{�`�U�k3����qD���RFQݦA����;AU��K���$@�S~�"�)�T`�v�R7�(fJ����� V�mץ�3ƾ���7�x�=�7��Sw��oZX�&ܮ[�M�c���/D��8�����Yi�ϑ�g2��,z@q$a�v+���0����%�[���^'�q�}��]h&�M\Ǉٺ�o�d_�Z��n�����(��iQa(-ëb��j� ����%\.E-��]^��
_�)�?�k0�_��u@�E���A�+=��B|�$�%c���6� ��/�� QPnG�ʢ�E_�� s �����kџY��><E��O����3d�v#:����0V�)� ��]���3�)�ep��!�:y�Z��s1����˳t -{�ڊu��Yɼ���E�����[�0�mQ��
B|yq��s�B=��BQ$Ƅ2@��ֱ�a��� �Y�f,��5��_��������h���R�]2��W�ޜ~����l�|�}�)�צ�"J�_b�J��
X��I~�Ƣ=t]_��ȟ�M�B�>�M�u��g�V�[FhPx��T� @�@Z���_���z�/`p�r�27-]�@wǬs4!Pxo��j[�������?�E|Y�MD3���j�U��aI�3��T轢�*��f��KzD>�����;*0�n��ׅ#����؊1=@���5��z�E� _�v�E�\�3�V�[.�H�a1�� i�ϲ3�x�����e�B�0�5B$	b4"K��Ncs�.��~�kw����:Kǅ�^쁰z~�p�Dt�H��Up�󀆲@�Z�H�.���"�S�t�������_v�u�l���c[����h幹�9������+- x�o^� ��9�68�^$�2nJ���=��K����v���<2�U�Yt���D�[�����fL�X��{������s�!��f��^3��a�����ά	���ld�6q"�~h͂1h�'�|Ҡ����c�Z�6U��2B ��Y��&�э�G�����j�yE�;O��D����q�0��!���̷�g:�5M��g,�&D��)m.jL�"�'�o���}�����m��j�(�^6&wh�� 4��^��j�|����n ���!S.�PFmX=�#���}B�����Q�}�Gg6�#�9l��@ߓK%�3ɸ"��;~"�uJx�-����p�
X=2�+����̳�Fp���8�$�Y�,IAs�F��n�q?�sa�02���<v�^BB�鏛�7n#�Ȉj|&�/B����b@|H@U�+X��l��˾`������.0�����Vt7{y��'}��_�4�D�
ۯ�N�S��V���裠�ݻv.{O �-�ege0�,,����=Q����`�5�d�L��i�L>�y`e�Z�u���}��:�q�u����y�JG�j�g�	�R�e�*��((�H�>�O*>Uj�G��i:ĩ�A�m����}ѳ+���w��n�.n��
\��'8OhM��̈́�Xk�4�A�s�U�$*3/�o���Z�
I�u���&M�=��E�F�t���ؔ&����j��BlH�dVԎZ�+�4���)�����/5�.�w�?Dp?S,�X0��GC#��=g4Dߴ�zC=�0�����g�t]_�&o��Dn�݄�pV^JecO�F��/g�ަ�+؝2<���*��z���˴�c6���a��A��[��q��)/S���׳v=�K`�/����r�pY�I�����;� �٣��;6yTsMm��=����N�`��Raέ&d
�`���f4�xHK{&�E�,fFj��8N,�	Ɍ��x�
3JM�F�E���4\��e"�ޟA�U�H�K�I��%v4ږ$]��-����� ��g�(��7�;��6	�K�$N�ѻ��������� %�>Ǟ�@x��=�e�bv��\���$p��B�s���@�"d|�� r�dT�`�&�7��a����=~hN��E��{�X�DˎͲ��r\�&rk` Q�G�W;fI'ڲWp���:�J�o�垩������+:�^~3[���R9�.z�}���-3���m�$��ȣ�"Re+Q�ːd#��seB"ɩ37μ!R�N�$�_�D�S�7�9����9ZҡƼ��_���NϝV��bo�oOf����=Yρ�
���C�|���Ǜ%��O�$��}Xf�P2C��/6����>�4���e��S�~�����,�� �z3���p��una3�"�Z4%�F�|C�����ÉFh5�
�����ޫ��''��|��,Տ���������y�G��4[l ��íG������V�gW���ij�X�ϝ��� Aˬ�լ����� Imk�lW?4���V�ŋ$c���*R:N�JY;=t0�`���܇�|$e�!�SupD�h��UF��X"L8�J;@w��_'l��S��Mk��q֗(�$Aѯ��0���[ EB��_ix��2��"O�^j�0e5QhKo篪B%ZE��h��e��̸��x[�\S��>µ�Q`�R��V �|��C* ,Ϝ�����j����"^�oo�֔Q�P��(官8���n�����u׈��L~�����el�ţ��j��'1�s܇k"�֗��`��-����^�\����1�ޥ�I�#	b�Ӛ0]��]ȳ0oØPRoh��狓S�բs� ��3Ij�8�Ɣf�`�� ��(⠟��L�2RR~t����3S#.7*flwY`�X��)��	�_�!kv��7.6�,� �8Lΐ5��T�j��}~�cDrI �X��E����F���jR<�:K��So�����s�$���R��!s,��I�*�su��b���{J�n�%�ԭ�'/"5��
�Svc��i��T�~%���`T-�A
�؃=��5b��ٵ�.��ײ�<�+z�v�^CD����iS�H��cRz�`��?.
ő����[�t��Q��0CHt��M«���O�����_HVJd��T�6��o=��,� +5T�c�&P���'���
�ī�Q}uYy��ם��g@U���I0A�
���p��(�`|��+ߤu7�޾)�q���ݸ�T.5���+�~�jk����[�����d���x�F���]�ʑ�@�1����|��$s]��6�g$��*\Ȉ��쵳�t��C�zh������d�B��,�6��R�[9�B���}�����q�g�<��
�e���Ԩ(��ݎ�G��r�Q�赂ȟ����V�@�[a1�$
r���e�D���"?p��¥'=�q̧�����G A{�?�煨:�h�ǯ�� 
)���7�`���0�:��2h��h��E�`լA�{�%��%�����ƃ���M
��Cf%s�#�"b�\�,�&�3���P�
m��2�Fs-�r���ܑB�A�π�S����O�?6�1� 9B�? $��b�N��y�R�)mM*gf�t�Dl�Lx)]aΨ<��?�$%���&�_:������ſ
)�J��Jh�5ʾ;�'�$��J폽���4���vݤ".�钄G�U������~;���&7�D��&��J-G��D��X��tC�<j5��AW��
��x�d�Қ�Q�ѫR�Y�ލ���� g apT03�3����%�����~��Ec�ۆ�c��1]�Ug�h\�����Wa�i"Q���jޒ%e�wn�X�x�>d�,�������0��[�v�������iŀ'=#��z|���z��R��B��I�zfDީ�HK���5Yk{�(�
uzP���x� "\*��Lq�nH�l�����Ǟ\C��|dU1|Q��M2�Dډ7f�q	���ăuL��hT|�9)�Gb�E�"N��,K"�E��>m�s�h)�(��������,�7���Ge���YG�ż��F���W$]m}N�d�C�G�iC\��r!�"!lCk'H j�/��v�Y�e��6+3��U�;=��釐C���C��Y���ȳ���/�dk]?�!�[/��a�h&�4C4ァ��o#$y��Ԣ�X�:ގ�p)0@�V㹤����(U�]5��؈���w0s	�EuS�\�B����e�]r"5cXe���'�Z<�/?�M��wy^ӹ�R�ʦ��Lk9n�:�M���ԋ8p�ڳ}L�DxD^\B�$M����6�1�Sv[���x��A4��Bm(e�q��V������+DlnZ*�,�Z{����>���w�2�Tm�-��,�/Fk��ga�.l�n�}\����Q�*��v���B:^W� hn4g�:�jaTU�h(ԇ7F�Ք�I�s�M�����e�1�y���a�F�W�~�|g%�/B���1��˲0�����>.Ǣ�%y��H>�5��4� ��!���!5L,�SO��{�����]v(L��Z�<���a�
�fc��,�Ń�	���ۍ��gr/�C�P�`Ooc��#�74m/�J�8M\�'����NԨ/�u���ʬ�LP�sR9�(P�~i `m�ݘ3P7�{ⓞ�����F����X�P�T�gYW�Nϝ�S��Yv�.S^���ť�
�ZP$&cϨ���*��`^=q��w���y��2�R=���"��65����P(qX��e�fs�ȸ2����4����6PS�E���9��;ˤu}�o�N��W�Z|F��d���gl��r�H|fʣ���P;�eB����e�չ���J���")9g�����w���	��4��9�7Q�E��V��\]�hk��
�.�� CW�WV*�8���j�<�m9�����%�ah n������)[^���q�����]��ĦF9c��k�s�㨗���v�g��~��g�wI"O���$]���:� �o�7���V��][�L]�ч��������$��Q�8��a���������6�2����%94w�ߗQ�'�J�;���Eʪ�ރH�����	I��a�G�@����b�L�b��9�j){{9ۇ��7�Q�G���>l��E�Ă�K�t��q�l�ÀQk����|��1�����օ_P��36nT"k��<6������>��6 �����)ݑ�Hz멎p�����*��H�%��&�(L�E���&[��$�["^c9`���>	�O��t��^땄�wI�J�����K��4�/��,d;�+��n�/�|���>�����W	CTS������&�&��ąRQ1I���)kZc<��V{L��F��C��ؖ��8I�Fզ�`'��T�W�|��~{+�Գߙ��Q�ݛJ�\���+�7@A�4��߃�b����I)�Z�9��4�$b>P��a1L*!���	�Ӛֵ���e��/��گz�`���1z�[{���F�	����l�i��ԟ���Z'E�uL�`������t�D��J,�.��8,R5�%b�s�Ƚ�D�]�K��D2�<m��F�^o0o 2%i('�bJ��o��42�����8.b��T
�����!*8�b�0̷��Z���$����C�uNX�A�Ul���?�u�3s��D�J�����l鼓^�c�ne�fZ���)κ2������H���W�� ���%�P}v*)?�:z�N���/��KG�z����ejĹ�ɳ�n�}�RMwx�p�����~.{�S�>���.�5!�/�-[��f)��_y�b\��Or�#�XI~��s��v`%T�u����zA�a���m������Lm42�e�ĈYΰsU��BB�&IS�K�'ǌ���r�����B��%Q�pl"�= �ǫ�s�����+�]�U`/z���#�Z����?z������=��WKp}M0�������aY�f�.�"���W6��6
�ru2������M,f��ܲ�}���bz