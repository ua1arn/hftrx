��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P����0��ܴ�t񢞦�Z)�7�{���O���Y d�7�.��I��8���c���׼��U��VѲY��=K ��#~q����4����Ĉj,)l,��ۅ03���c'b��#I�Q�K4��KB. ����u%�7�}�eTB ^�����������W�|�1c�*�K��g�Zx�+c�_9�&��O�1O�Vج�#�o��^{���2��X��B+ӻ�i��w�
m��>�麖נ�^#�"�
o�VI&���l����~�B{[��$'Ҭc��Ό�̃2���[���<]�H�@���ɾJaVh�Z.�v�el}�(����@�a3�v~NO>̩���i���QO5�gR�}5�$>~��!�PC{�<�!�"��s4�\Usy]Z�c荱������>};��h'�R�ճN#%�O7����f���k��a�*y�Y��[D|����#��r0�j��U.�!�k�,a#�N2��@Jmi��^\G�[�V�5��<:��,�e@m�/�F���ʿ[���;,�KDz�N}��u�H�3�K��W%-�ܸ�'�~�ޗ�Qk��w�e�K�5��Y���5<��'}�)���(\��{����1�%�"%���GZ^�U_Z����ZB��ؚ|�hd`�xƑ���,[�ClyW��U�.�#�4�~0�0CGU(� ��Y��D	��/�z��_�AQ���y?���X��� w@B/��A. ����Km�ȺkC��<��}Ű�b��]E{]���[9�i+a��|��R��$j׳Gk#fXuh�**�wNԳ���h��*;�iFB��	 <�g8���WE&h~��d�Fs'�yۗTD�>_~3<l�.pR����\�����v-�@�c�t�QF�ۑ������q��y&� 
P��o�(o��5��c�2�1��	�OP潑��O�jIF�X�Z�o����8!Y���>k.,�=Z�_���X�}�4�1�kfr��}xn2�<6d��W�Ш�Oz��ˮ����F��x&nؔ�Z紹�ʫ���s����ݨcY�oQ��!�}H�g�Qq������pMxOI�j��&NЀT6A�
�?OO���=��N)�A�h���SQC1����������*b���YF�!�-oI�Inm$M��MnFi�0�?TР��ؼ�Jm���@�)�L]�.�b�|�|
s^�?^��!��swX�դ���UU����GiQBg�M�����z��E�L���Æ#������M�B�Sp�\ITQ��|<X�����_�����و����o�\��8'�F��R��9�Baǲ��Bk�W�IC6W*�]��ގ�Q�`q��䔣�,	�^�YZ�c����g���*�c��;�����o�H�*@�H�Y#�����%����-� ��I:��%��>4j��.h�n�Yz��)�]�]\��f�Mj��fW��T�s̵
$esj���Q΢�ĺ�`` 2s�)�b��5=t�\��,���4�/&�RYs:��ĨLFR=���O9_Ix5
�0�n|��#�|�ûA�\Y����vÕ�qC�#����"V�:�=�Qk6�э9V���|��Sa �9�$qR��a-�h����X4ĝ+�C��Ѱ"�w�;Dv<����l���C�}���S�̠:pt�p.�T����j�u&�h���F4+�B����Yoa�Tg���G��NPw9M�!��M� d�z���s ���04��'�R�j���G�-:-�vr$P�Д���7h*�n$��Cťk�e�ǕrכH�*�>+�=,,4�Og�GN��~�����v74�b4F.0��p6��$/����0�R0� �6!xm�8'a�D+\�LRPe��2�#7��+���5��� ��N���n�@�t�Z�\�s�9:�w���Y'{BZ�k\nR�77+Ut3���yX@7p+f&0(�Y����d���}$V*Ը��y�WՓ��2��_���0
�%��9�{x��?�m�X��J��H��ع�@o]�Ԩc�ᛞ�c�����0���|���ϧ�4�d�a��
��@S��l��o��Ë�M�l�N�	0�?(=�v��3N�o'	������h.��Qg�65(����1֋kcڌ�D��ftv*j�7K��S��l��_kscǭf�n\�����ai�9>�<�PcҠ���w;7�@r(y��F�<2���m�2h���}B*�j_��e��1-Ú�`\נ= ��_����Ҟf�E=�d4�I�E��y ��m�*k@�"�c�v�Q�Ǔ�E�R�HCd6}wF�d�0�]mz�����j�o�j	 (�Rq|�
�O�jMۜ�Kr�OF*r �X�~U���J���I�wq�Z�*�zp[Q��*�(F����vh.�;FsrvA�rkF���x�����{�:?�0�s��_b~�����W�E]��� H�gڍ[��}���v���k��\���	}��r�,�9��R��4�Dh�����u�_�L��@~�~�HS���Qrס�z]��=9s��g�"��L� ��ylݱh��C���zO�^���zB�R�
�%��0$R#�����^J�:`jeF��o��rY\��ϒ���S�E��JvD��Rr[Ī�T�h�1��bv��^��N���j�\G��<H�_�}���Ԫ�Xyt]�{��yk��B:l��R����U��{�'��ɾ]D�'���2d�'ǹXD�9���j��?�>�2���

lu� kb�b�y�#�U��Ԋ��g3�-�w\�b��n��žƒ�%�8���a�0�`������Z#%�sNX���6����m �B�V��&�(z��E�	2QL��ek)��?���<e��zݹv&�LUk���2q1��\盲��I��rH�,�̕��RӚ��;�t��%�؆���W=%c�˚9����;_㳻w�輾 -�<�lRH�k�S�C���G.���Q��]� =|Z{��c�pˤv����D�^��h��c3w.��S�/��$^�9�|G+��X"��2���}�H�p	C�A�(�LN|Xݻ^����N�D�F ��Թ�y�h�h�Ш1�K���X#�2���1�I���g���K�_�9p�"bܓT���9�Q�+����i5����h�c�*�T�x�0A����� ���b|k�S��C���lh#���-!�ͨ�|_s�Dx��8�Z�ps4������,t7lP?\��tp�$�jy��P����*"	 ���"7�x��K�I����s��T�q0��R7���]�Ysa�����)1b�A7��@�'ַ��q�c0+~[�1��ұ���(�8@a�"j"E����K��j^��J��֤�;eRø*Y���Q�^���P*��?��)����\@��/��ӵ�a��|��*S:N㫗%�n]+1��.[Ni:Ҍ���dl"?x����pI%�� �e1O�G�@p�������ӅI�벁�&D�eg��K|F�4��\��Z�Z�(�����Y��c�m���3c��n�Ss�^����g����չ�0�JΨRE��82���}��;�@e�\�l	�jN-Xg(3tSEp�(�Y�G���K�W��Θ��		��N�4���sA�A<1=�����p�f}�o��<n2S�{x�ܽ�S���s��;u.�k�AϟW�+��k��`��Y[
�cF{����H�hA[	�n&֔l����� #䇢�/�7�o�6+{V$_f����~}Ak���4����+�Hڻ�X�sMD�BcF�Ymv1���L�|���<n��o����8E�>�x3���kr�S���-)~��R�	6Ϣ�em��@�:$!��P0�).5a�s��?�0�3��Y�W��(��T7�f�̦�WѲ}�=��Q}.�^�%ֽ�#��S�+I٫�w�i��O�����[s6\t�,�M�K��Dqv�Wm	\3w覓��O�; ڋ�SO�
����2Q���"�ٿ�_���A�r���So
R��l�JQ0'8
��QL��k���g@Ke�>!�$aAF�FIiT\$.�*���Y俦H��?��W��3��i+�֡�.ռn��A���(q$^��c��w��K�X��zm�gK)��>�̅~�a��{:�hH�
���͔P�s�*"�z�a�c��>�
��eV�}{佑�X��	*W��
��!A���%�m�u�����F�IK��~��2����OOv�d���ǓL
*���ٵ�ٯÖ`�Nֺy~O�[XQ���Fy����]�n�Ӝc٬�!Y���v�2ڂ�x@��:�.b-�Y(�먅�RE]�1]�"� ��H�Ƒ�x3S��l�샿�*ȍF�ci��{�u"Ϋ��f"���3���4�w��3uH��PRn���AY��|I�w����O����&����7��y$��������#;�Z�r�C�E��\*�X�^�£���_یP�f�(�p��L�c{Իie�om$�k��ߡ�xq!��L,�DXՇ�s�8�@�#1F����A�R���l�u_�[:������"�xS,�h�0���v�*v�%e��s���NeYP2E�.Ą�C{��)���Z� $��_��~p}��C�e���Wp-*�17�~�'����C ZuYL������T��O�"�b�6K��G*
r�/3`ߞ��?�M 1�C�q��%�?4ć� ��7� �w����,�\���ni�*��1�����W���0��x*nNr!���n�f��})K!�`&�����_�p�?��]Bt�at2��V�Z�d���"$yI3����GZ��A[�i��!�-b��{��H]�-�3�ˈr�tw0��7��2���ͥ����'�8�0���&qIU[��#�I7%I̐HJq��#�C��:�TL�r�	�
�'�r��s^��"Jvja�EӾ�M��� ���̳�4��Ҏ�9���x)�1�����b+��O���7�+Ȼ��1o�+�>���6����JU*�R6�J�%� ,���OP!~��b%�񐪩�/lh+��	�-6�9�T.��Q�����y�N e��,��|�ˁ�7TB�@C@#�YH����Albu� ,F\I�����~��.r<	6B� �],h���ّ�TҖ���8����]���M"�5C�����K`٨~^�����!�,~\r-����*\��Ϟ�s���*n
�s�L\-s����Y;LW��}��Ȓ��!����n�:7�E� �a���SM|�����״�k�!Ɲ*M�@�p���ѫ���O>7dfڒ�8&�b��_C�Y�K�S���m��&IâdꝆU��d��}�-}U;��`W5�HEBƯOa�D�<E�����l�Ec��f����Q��C�[�=F3�%��l�D�� �9�J�PWA¥�������?�rH��h�J�da3�a�6�C���G��]���n�ɦ��EC O�)޾K�[X�T(��\
m���UW���%%����#�$Rϝ@�$�"��#����r���2V�N�"d9^��D��bN_����>�Xk.�"�!O�	Y7�DG`<�AK���ʞ�Ҩ���������.y�.ݺĠ��!Q��bB�^Y�i]����gB ���J��T����sn��>�͌"����3<f����`.���b3̻��=%\q���jL�RV���`�@f�UC� ^ـ�ǲr6�MP��L(����ɍ����tn�Ű��J��ͫ��eqp3�S�Wv�e��^���(��х����a~�X?�7/�9��i�?��b��.�l_��^͐�׾���M6u�lƯcl�j� ��!J�˒m�?_����=�|�X���	J�NG������Ȩ�ˏ
�)nˠ��9�.5eE�6��y�%M�	+�^���}�����K���*���} e? �f��2;]n�
NSb�]W���H����4����d�V��ٯ�(�g-����V�3n���3 C9$~sRZ?6�Z
Ĵ#�J��w��華w���O�B����]���Y��P�� �z/�-����o�����L_t�����O�=E��hN�-����i�m�OO��j�u ^���x�>�eb�ee�>,�}��:�={H)4��
?�!��?��ݷ�w�-V��lj��L:��㸤f�4�����x������h/��,��/���7�Z����A9�/9��^�; X��TR	��Y/uQ���|\���s�An�������y�3~��>`��߮�d Q�x�%_��#�Q��V�e5�1����'��Y���f�����^4y��{1pUq�|��t����AZy�2�v]���p	�ƈo��;=��D�!cw�U,�]D����<�S@��