��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�b.�B*��]Q���n��4��$�bJ�3�`R۬�U�-���fMμ�al�{�"|y���.�D�T�H�H��U�J���sR?x�V溟i�+U>!㶇�}oC�n�����3�>~��a����Y޶�G�BW������BR���3�v�8�y�Fj�,�8<�Cc(�(���,��k(g #֔M�!�7�����%OC�_������ا	/k�Tw=]�m�B��͏M���c��yC�uL����+@����;�S��˅�*Z��]�n��uz��V�ڛuw�+S�j.�؇�l		0�6��ZA�nR&��Y2����;mI�L�qU�7Q��Nl���5V@��)nI%!nΫ�)��6�i�`$}ԩ�^CV���E�b֝xr�=�$Y>�d)���l�����L�g��t<�4�}��ٯQ�a�;�]������vW�s�Y`� �P��RGټ�
(V|B��]��p��ΦMXw�n9֬}R@:�*x�VX��+
���W��\p�ک����#ĖJ��1X	�nH.���;��0_�^п�l����������c	t�o�5q�EJ�?��ҕ�wI}3x�pn��*��¤M��	����	/Xl6fh�͔����~}t6���UL�Ѫ'�e� �{�����H�+$�8����c��AԄ�\x�!lx�%��͎c;�6����A�4Y�.�<�w�c�ݗ�X
	p�����6"[,��١��y���Д��&J�E��1�\/�f�����t�"@�nθw{5)>��*���SM�ȏ
����e���A��H#P�G�c��_���04'�0��8���mv�Ƣv%; ���eF���5*��������2x��|hǥ,���R�Zn�s��,����WJ�obX�@ ��"0��}37����G���٭�~�%�[���r4Iѽ�ܴ����j]y�_����#�IL��O<qO�q�'����|I��C���O�h����o�Ƣ������%�> l;f}v��>��nTTX����u����� �к/(_ѕ������ �%�65�kY�-���[ D&f�_Z�$�,L�׻���.��uv�j��L@�=�S �¾3�P�ͤI��#��V����&�`��Q�orƵv��KՋ�I����AG %"���8����p�\G��`�`��Z�Ֆ���wq���kp�t�IhL�1��ٷ����8�p���/���N�~�gx���qb��v�6�0�6>
���k�.�AC�Ñ�'�4�ޖt�����~
�ƌ%� ��߫Gt��L]%\�>��K^�;90EU9��R���`r'W���8�W05䣩�W�|#�XZBf�(�ff��0W8}��|s����I�Qi� Hu���«s����qi�K��E�&����}e��?N�����U����>1a�<u��Շ�҅��KcL.�}�����Ve�ݢ�EG��1�.+�}
�t�4�vb�ƭ֧�]�t��1�&���4Xf!1S��W��=�=v���@�<4����9G?�>�䠯}}��Ӑ�x��jMC�wS��GFb|Z�M-|�*��
���zrer�Ʉ����v���	��Ο�����*���<j�F�fѧ�S�����%��IF3!�j���Ɇ'+��m	)U�t~�9�����<X�я�Ba�+�R
�9�9�v�����hi�ID�mY�CL~�%���yM�Rv��O���C
k�C��S,�<����+��$?���P�Q�����e��,݅�e�����j��k�@k�>y�-,;]���[X��$ct�n]f���֡�2��~��#�W�Q��I뭓K+��UG����(6v/��'b��N��֜�Ogk�-�h��3��vⲋ�ؘ9�O�������^��e	�t~�-%�Y��n�JU��=v�3�{(�ih3��4�<(o��F�$�f��d5h���7o'�:A�Vo|������%@�$s�(>���!]� �Bd�� ���xGs��](hK��q.;�=���!G݊����m��;����\� �[wh��[YG�k�Mo[	J2F�ϐ,���{�®��'��3?{��J�&�D�L�l�]4�L<u��0�}}\%V���_`e��͢���~��TJO�4wB����-:_�g�� ��~��i�ZT��3S&"ɂ��m�����;��%�o���2x?
zHL��̢�Qz��W��an�aA�S��a�e����:�m��n72��t��ri����
�×^֛U�ݖ���g�	D�M���R�O��sѼ͒�v���e����exј�e6
#e�X@*|�t<B'[�_�i����7�>ڧ��h���?7����&�d���1�BX,8LصZ��F��(�}[>�kU��^&u��I�[5�?�ub�o:���j���1W�{�SGl�S!P���d�s�w������ǥ��J*��g/A��u���� k��yC����e �R�� "{�"Ɯ�舅���ӛڞ�y*{�Ս���W�j)�11:BqL�E��n�
p��>�e'<�ܱMm�0��L/Ke<� �d�ߔ��yzo�HD|c~�|]FYxa���]V�gT���7D�Oܽ�8��d;�ڶx8���ۖ��;g,O�{`I�#�ۧ�o��z�pR��������Q�t\�U�INmB�SF���yHU�{u�'ɗ>��@9�r5����Ea��&��@�;nS�l�Pc�6<X�X�Y�PK�D�#��fw�AW�p�9J��gH��.߈g��)���;T�9�;8�I4Gj� ���2�*�@���ʐ��������A�i�M>ޒp 0m_4�j{��R��p��vM�%��2�XT���o	m�0��/'�=>����?�R̓�w(�&^F�B���G`#�<�K�X-G�{P�:B����D�5L�F�/S��8#��(7���'*ؚ氍�P��?�dPb�O��Fq��oE55����
��P��upGvvS�h� {Z���
����<o�*w�r�{��%j����l��֥**n���ך�c8�z9%�o��h���ƞ�u��?u�V���;"���l����V�ĪTLH�EG��񤐴ѡ-s�!X}��L[@��<Bő"�0n�k���#�c.G��]H����8ml�8��өY�]ϕ�>H�91�W-	�f*dMw}�t�]D�?kQ��2l��*튫�����Yܚ��r"y0�L���4��\L�c=t8��
�E��t��d���x�v��by��.���-	�N�g��F\�(0�J��$���Bp����Ի��u�Z�:?���p&*mNx�y�b���.[?OQ�� �3�P�צ%�y�h��g�X=԰w,�PQ����TGۮ2W�E��N�:gwK^I���߰8u_9�Fh`ۤ9�#�<Da����6+�`~t�EX^>����EQ��N�DMJU��knו���=����]e�b���g�1:a16��?dt,�����i#�����M��wR��g�B����A���B���Bf5��7)y�{2A,QY��do�_,�͚�>j�Ө�Lv�z3Da�;��R����H�ƛ�R^4=$H�7t�I{Cc�l���P�,	zh1cH/c��D�ר?�ڬ�GC ��#���hLC�B̺������L��[*
K+��d�0q3��6�%}Se��[��� ��v��Ql m�7*���
�L̈́�����H���g655V�y���x���
���Ps0m3~�7���4Ґ@�ySy�����=.���c~���i�:�� ��6�W�H�;3gJ;���TfI�VbkpE
���T���T���b����"���̌�o .�D����"$���,I�@-��
��� �DDP!��&�V�C*'���"���v���j�T�̸�`i����9�H���TT�����OZ�n^D?'!0@5d��񿍂I%��}UVT��[�Ljn���Fk��0�x8�(�A4G+��C�L 97o�I����9��8�̨~���%^r,D�/x/������c��t��zA��[=|JE��`�R��,�Ҹ�Mc��g�6��l ����}<��Ņ� �:�-`�}*�1�u��r0�+s#�I�}k˕���}����Z��HL�iS݉c�~�
uy�w]['����z�N2��ǟK���5;^T2���y��Ē/y���tZhY>�_8}�Zjp/9��o��~����eNh!���W�\�&h�W�P���t��X�� ��% �V<l�+�H]����Y��@'�fѤ������p]��E2�Eo��̛�{�S�S���8��yQʜ�mp�a�k��-�E�O��.VQm$֨6���2��"#^�;��,�懺HZ4��_�Y�S��ެ� ����ȗ�������*z�1\�n�$@b{Q ޞ�0$o�C}�y�{�c��w#f��R��.ؘ%;�Z��C�ҝz.*�5 �K:��/j��$�J�RևW�yq�?����[Ӛ�7*]Y�������˵=��F�y�$�2���D�Q�Z�"�>��l��xz� �hY��c~�:���5�C՜CP�\�A�M���7���0���rf���'���m���?7a5.�&Y�HbѽA��/t3��O"ް����d�ĭ�H>�Aς��}�n���&�V�ZD=Uݥ�1��qVC�k�36-�z�S�#���Qr+\

��E>�n��*U�&�[��t��.r��Q� �fJ(���K��Ε�u@�#�vCX�B���m+/˰�U'6�t�����b� ���Lc�\��(*���AS:2�� �g�uy2/ja�F���ɯ-T�]��9ɧ#0�?���+G��Z��(���{���J��$��m酏Ҽ���XJ��s���Y$8��i)��s|pn0�%�#�Bn��x�H_��h�nTT�M-�Q����X�d�b�u�aT����G�N`Z��C�h��ä�k��* �>|�[��H���{�-,�Ҝ8T���螼Y"j����BFܸm��J=#-�ˈю��X!�~p��$�i��4;�09�{�������-���ͤ2e�X�77��]�����#u�-���p���"�w*0���VW�s���Fv��j~��I��q�����Kf�s������e�9�g�����P���16�;��>��<;�9�%D���kh4����޷?�C�r
D�)5�N-]n#!`��W�(:$�fY�(�Y)J��?e3��^��%�j����Zل�/~2���B��mő��� �<�Z���2�7B^<�Dύ7����c��l�
%��ث-�)Wk6���
4�M��/n�'�/�}J�]�PO��%���q�B��k�g��2m4��stsi̡�D�L��X������"��y(��⽢_��̾0��E�2�I�=��˗���+���O�u���R�J���;_����Fo��h_|��.�3j�ݐ]�!�0�+C�p�VY��oFn����Ώ�ٹ	�PՙGP��r�DlD�5X�U��,�)�[�,ڡwø9��wKt���"�\*7�Rj��%W�
`b��|�$�c���aϖ���쉒I!81	7�s��|@Q�|���`A\quĥfS+8mŐ#��o������y��E2��8��kd�c~q���wC�}��	�i5��h��EY0�������=X#��a����M��ϫ�#�<X������f=��3�}ՉU����V�N��Wd�%�C�H��cה"ZM9ؚ+�!��T=kDG���N' Q17¶i6'�v��?c�< \�(��zcJA��۲���wQ���8���k'g�b���&ϚN�!��l���.���i��9Nv�D�ib[������XL](5Aȃ���$�83���[9c�:QnW�r�vdV�	O��mճ��
�/����T�{Y^b�x�yd�*s� gCv�Q)�S˪���Y*�q�N���i��j9��0x�1�J�l�'�cWN� Y�f1��i�ѿ�{�3�+=�3'��2��@*�tZ_0���=��KӤ������<��/��b�[�����`�8��	���x�̄�:ak��Ha�f��n.Ķ�n�m�?5��CxU�G�N�x��k�X���*%z�;��)�#�D�ܜ��B����-�9���Y�膺� mY�2)CC�E�5���#��ڹ?�ZA�;U����ș����G&.θ���xi��k�����%��E���������^@J��-��({�I��ָ��H��ly��t��s|���ss2PP6 ��~��ձ��i?pe]&O-��G�O8�f/�~m5fo�����>����	�8&�y�Ss��{�KVD�|+�Ͽ}��l�4��Ux�Lg�63�}��I���-��S�T���n���B����1 �Ui
�a�9(����}���Y�0>P"衖~�qUB%r#n3����$_��w���n)Y>��Y6M}�(_g]������)�{gt+(�2��fd���u4_�.
�\p�W[� ����`�svR��r�)�՜��4����T����л�W2����>�3� �lpi��l q}=�^`+�4�i	_����)��ש���~�e���\~�|���Q������}���~A�~o���|�g�$��h+�(
q����w��Z���x+��QGǟ��[�%Z���Hk�5��9t�a(Xh���Z���)T6=X�ٍ#LK�竩g��)���+}P�U�����ǇPWyt�3H�c�O�ƾ>I��Ɓ�Nm(]���ӔB�;*��&����!g{C�:t�́4V���ye�T�a1��Ϲ���ZӃxo��;�!*vQfp�����O6RX4����ś��ĭl�!��>6��n��6X;q>��l�>��Vpuh����=J1���3I��6�ؗu6���[�,�ŚG�#;YA���Cכ��8A:�
~���EG��P�T�=EC�k(�#H��3K[n<�9a�㞻s㩮�ӆpR�3}�*{�$�*���)0��e�+����X�����u�9B&�L����" \"E6�U"b�]-2�e������ L]n��R�W��/��I'���Y\�Q��KE~�����2L�6,��rs�����q���lګ,*�8�2��,�f¯%Z��Za"�+�'R.\��~`�"C z���hM��ek.��I~��� )�y�S,��h�x� ��s��ʢl4+d�IH<��A7��\籭x�CQ�ƣ?�{k��#G��d�&[=A��`\�\��Pwn�3[ #@���Yk\�g��`���6/�����|V̚Nҳ�7�r�"̐D���ܱ#"����4����r�����؝k�����<��4d�-�Yk���'��-��d�y]D�"��
闣�EB��>(�ϪY.�r�%��f�*�Có45�R��Dw��|��O��($#m�@&� ��`�N>�1]�avN���ڢ7�y��$;7H?��0�F��
�����@�je}ZW-K4���!�v�B��{�d�;��Y��Q��+DL��J˓�@e1A����~�L!aۉ���F/em]�����!���N�*�I��������;��-���LG�i�^����cf"�}�K�	
�����g	�ODQ�-�2G���j����U��@��f��}~��*���u]o"D�}8@DƧ�@l�A��;�q��q����r��¤�`Մ��E��1X$���B_)y}e5����H�Z����	��U�1X�3D![���g5�]�d���rc��u�A=�|���ӊ�ԮJr� 93����N���-�4ؑ�Ր)����+�ЕYM{��T*���u��I���s�|���}�U��p~� ��n��ˣ��\h�j���+J9��]�t#���m9�h���Σ���LE//s��I���Y�Db�(�gA�ɒ�a�)Y����ډx>�"z�x4�
)�y��� ���y���0��f�Λ�P���!��������Y�b;hZĘ^"ml��k�%7p�K�qE8�[ t�3�%�ák�ù���N�u ���<Ld�0]'�GYf�+D:�C/���&����(&D�w�Ǖ�ٴ VsL��w��ļi�_!b�X��Y(�Tҁ�,0�g���i�Ko��ڜz\e~B��>�C*)J=�uM�7%���1Ec��@������X����YkA�� �sHoR%��}�v4���Z�t���rr���YO�yA ��;XaA2���:���V����ie0�V��~i��>���'��@҅*���;Ȋ�V�����x[�(/w�d���'Hke��uD�ҡ[޲�Ճ�q1Q�����x��Z��aDE<������}S�9N�c^��v��K�4�.+l|��~�inB>k:�?6W�B��Q�S�F�b��*��$0u:#d��Z͝{��Vx,U����*�6ENj���M�G�uU�Ps����W���i�T�C��ʀJF3YX��m	9���! W󎊗�ߘ-�t#�S+�8zPF�&M�M���hd�F��=y�#�a��E@'h�;���2� w?@W/f����^��W�E�h���
�����W;�+Ԕ��1X�	�H�%��!`����62Ȉ�����/֝���a�١���́����0���w�ő��)���3�	�)�`�{-@&�Z˯����.9OT$i��i��	�
�ܕ%�P�E��*eB��>,��;�l�Ra�j���u�|0T�����h��� ��2M�?H,%��,LX�"��ڒwa9�8,�qɈ�^]�na�r�x߃����n�,���&��*�B��NW��}gb�2s�AD.��c�Qz�r̈�PS	�*7H3�����RR��ԑ�ĕ&�l �o�R�9�������h���?V4��q�k�i�̘Q�oԿ��_҈�ֹ:�%��s9����ΗX�&ް�FƼ�X�6(/�1F���[$��Û%.̬�܂>���]{4�˨v�����씒�����@�=z��p��O��.� ����('L�dZ�����/�j�-S��S��Y��pD�~����Η<�o�2���ݟ�9�(O�hF��c��	]ki��1(J晴����f��f��� ��C	Bz4k
�jw�Ɣ�gW��XG�`*y��9�*�F���W���}c��k��D���rFf�G��ʊ 
�������F�Q��-�̶��`[Ed��g�!��D'��n?�O-�2�C�|�J�YW),7�d�oNb�;�e�I��`�BԽ���oj�_I���ե�\g 7�'��V;�"�����|��=�w�Ugi�6�����u����kp�jf�p��_Q_C�Z �+'�H��%�?��keh�
�Wi����,6N{ˆ[vK�MBCA߆���M�e��M�/,>�-P�~�݃��m^f�l5sH��oڴ�4�ӥp(G�^.�-;����͊�4Rx[�PQ�=}�1r����>�P`��0�İ!�4������D���M�dN��ӱ@Q��m��n�_J�"���n
�R���6��4p����g[O#������p�	�TO�M��M�j���f��j�飰F���3��d:�bj��HØh�΋*"�Nf��!��|p:G�羠�E4Km
�w?����d��H�l�Ͳiah�<u�X;d����6�Q�tѼ+���J�n>�5�����$L��0���C���@� #:P�P�	�_� m\qR��ˉ,D��[,G������u4j���CU��A?��/��uv��6�y��+8՝׿�����K�&TN$b�����q��)E_�7|�dE=��a��[���9�HƪePf����,�'u$�
(�o��R�M]g����خY����KF���t���6MÌw��o��	h`
�ߗXC
PV:�j��K���x�LN�ߠwF1Q2�aya��se�vC���h�w��������[��6�Y?P�O�~S\Ҡg�n�L���������C<^�4�jk� >����f�G�\�DUw�%�u�����k"YjZ�p fS���*�7�xe�hs��
�c�N��|z_�3�	58�"������'>���Zp�2P{G��<�c��y�{<��b�^Rbꖥ��.K"�]���6Psg�h��.r���L�q��BǺ���-$KՊ���.冟�儡
:����W4AGG^�B�Y1ٞ��؄w���k��7�p*^�
�֯,����L]�����`q�&�}���j�ޜU���y�����h�I�l��jMN�D��\������6����ܶhE����;�R[�l��Ⱥ�T ����R#���������l��; /��]�l��lH8����:�'��Q�u�n�� ��s��_�ϐ~na�E�V��o"�6��)ם�a�CH�Wv�2�6 %�l�C��k��d� G~n�ꏾQ�����/���,V"J	�1 �'~�ʉ�D�<����1��r�.�aT�p*T�v�T���7H��C��F/��{� ��g��~�&�W���d��ߎ
�Q�%F��ZBt�(Iu�s�K*W�@���詚���N���>��l��ś��t3xT�|��ӯ��&W1�@�:�M�W �<��-�)1�;{ 
�B�G� $Ԕ5�p��!Fd��c�WI*����̀�z�59%XhH߮=��ж����a�+����V>Uy�-(1T)f���g���xxq�x[Ц�m����:�)jh[��0��,2.Bݑ������\W��Kf}*�b:���^P%6r8�R�}���	0���T�M�KX_қ�گ䒕J@u�� v(��)�>_?�T�u�?Dr�z`��$DJ�Ys��P�"k]��&�5�#8p!$4��u��-�z��������©��XsL��-�T�����R%�Q�2(�9b� 3����kL���X�~�	コ�H
�?�@���3C}�,AK�o�#p����T�{;��>T]f�T憔"mͶ�5��=��k�C=�p.�����ڑ]M���,sl��HB!�D
���b*x1@���	�����+Oa��8�B�mVd��b�0��6���j��л��ʼ�E}zcYpx@����;��Xİ ���H /���������$���\^� 컍���LM9�]"V�#Uo�l�n �{������(�y��~����s������t2n�Y����Gm>�Q���d㢮���_6	�`�Sʛ�Aٙ=��S�T�\2~E7�ADe��3ݧs\���,)怷��v��=���zGvmi5w��ʢ�䐛*o��J ��j���9oBϲ���:��f����LF��Zn�!|�Q�UMQx���Wo�&������W��g����{�5^��І�5qqp��}��;��}˧�o#����F��dT	�m��[��+�*::$Q��>Rx'��]ˢ�fEа�[��ޖ���CW�
Ӕ6��t�"�ӀS���~�s�$s�vM�%ʏ彥Q�ŋ�����(���{�;�p�g�oǪ0���#&��Ψ���A��M�q-�ײ����0�Po8H�����Z��݄pLHWo5�`��N��}�	��յ$t�p�T@�>�ҰGdy4j6a���=�I��M��&�E?3�2�=z�W�L����������&<��4�#�_��ˢT@\� Z�`�up�Qu���{����2(���a� �[w,�߼Y&1�\�lđ�5�����?]B��'��E�S�p�;V��VA	�0eַ	U�#�M>/?�~�Q�-�!�#�Ǥ��j+W/�4��r���$^?%�>�����s��	�:+�Kfmt�,��r��uHMY��O��Ә��Y6G�����.��(0qG�!+�r���mƥ�՗��qE�L��;�R� ă�k�H�f\Wuu���3�=�k����h)m�[��������'�'�i���Z���"y�:�a`��_�Ժ<N�� �M�C�,�%K�����G���G�`��"ǫ����=��h���8�y��e;(T�� �r���`n߮��x޼��x�
+«��ؖ �1�Gg1��-e&`��"����a_�њ��1Rx��'Q��P�`�1z�K��(ZL!TЕ�'a����j�\ίG�P��bfoB�z������l��!��(OYu�Mv��H��-H�<��~�[D�"Km�WC��oNn1,۬Po��i-f<-��#��}uuv�����pg��e��UY{:�t���%�>�	���m�-����[f����&P�CwS��W��d���IkS=_��_�]J��7�Y���G{�d<m�G�,<K9Fz��w�RHw׬��|eB��V�Y,dc�_5����
r��D(�6���d�[>`�q�,`�GTQ�	�߂1m��
��Rug'k*bT����B7�'�Ɍ�n��ʛ��]gj��HN'cQŌ�5�O�e_@���<�y~B
����;W��5���>l��i>=#(]�Y��11r.䈮vB�7:�&���".췬-��=; �96��������A�)�9����Ӊ���k�5ޣK�-�'gq���ҥ
�pA�Ґ\i�$Z��N*�kD�5���"�C,t�e�މ�G][=�έ<H���!pˣ�t�%N==�!��T���+�Y��sa	D}�N2F@L,\c�Z���W���ceU��o���bBa���ځ{���y��HQe~�,2�(�_s��)����wX@q��:����w&;��*��p��	q�+�)@]
H ���K��:0�m��qTZ����`	f`-�}�ڃZS΀��!�C��=���2��arH���7m��3K
a
Ͷ�J6�uAi�D������u9����\��&�S������m�'
K5~{bt�F�ʿu����'�U�5#~��]��ܘ �x�0k���϶*�iLu�'D9���yʔ��Sz5���J�=T8,¯�$�&�����%�Y"	y�
:�;ܭ���Ec�Db��%��8�;Jbح*�Y+��t{n�K� �BkvKva�Uٕ���2N�[������r�7�����t �>��w��(=�H�����e�m�-!��<`}~�)���M���,�X��^���\���o�2?C�9fǇ��.����kɴOq�D}�ǄC꿣&Ha�0)2��N�T�M��2=}��ܾ��&�����Y�m1��\W���J����d.��^q.-���A|�2�s��o�`�/q������$.�<��5�2�}8�C��1���L��&��=e#�YBػ ��%ͫ8�\`��Wחc�X6��5#�!��A��WTk��&�vr�|S�ٽh���S:��/�$�Rr����K�oj�bc��3��}M-��TM�6~�/Ъ[Xʸ��x�����o5��עl��DM��wF��p`�F��U4�mofc�w� �f�*�/:K�'C����,��\n�2���pk#�H1� ��1p�hSNܜ�|��:���"��L�����='�fLBIG+p|�D�fg
�Ҏ�]�`ܸch�z��6��_�s՘7�au�H�v?�ď�QE��A����Cy$��K��/���v۽dT�@{�����Ń��Xi�R̞#�3�9�?P�:<H�Ҿ���7�9ǽ ��J�)1���8�,J#v�e@����:p�SZ1B�`�&K爑�ứ*>�4�'@��V�q�¹��@��B\�\pPM�zG��bh����:Wlԧ��ix��?��R��v�ʠ��w�,q��eƘ5�z@�ߎm�<�w���4�f���n�[���f�jR����z5$�V:�e�8��񪹻���>��f3sB<B�M�YΏ�"�����|���w[pNy������#��{q�/���
%��E�-1T��>̊f^����&k��]zmdl�2{0��a _i]j��I3�Y�Tใ�6��|�׆6]-���v cUO$��{��`��q>H>S�ϒc'u<o�b4��ѐ�Go�s����I⻤���U�agOQo"e5)sB�í���>mȅ7���~����\t�W=Z�ҝ�A�>�m��>�$PU�~$�o�J��v�0DL�l�U'#��C�N��5��%=�4��v�۬3X:�#�V��dP˂UꩃoÒh��#�Q\d�� Sx�n�Q�Ѷ�������S��v�{��A�·�i��jl�ˮm��-R[�E	�]�����zHK�h�cZ�){��5�ds܇��۲/v"��l��8���E�_��4D�U�k X*
GyM�8�*ZN����>���rｬ�}\�ZM�������&�I��0��6.o��h����0�4��v�49��0�����b����g���(AsyC��F��H=���jf31x�f'4�@��$�6�+3A���I�y�n~��$�r�u$o@-o8���:�����	�֙���5E�IcGa��f�
{bؚmk5��7"�Ǭ[(ۙ(�:o�ڴz�~�C��Uy4��n��~�"k�.7�3��6��+�� un�#�b�o�H�=��A���G�C�-�z8ELjGtQ=�DG��O�פ��5>4���<b3��v������c�Tr��Q�+�?����2�[7t�33�W0�09�Cה;ʋ���)�Ηm`]�A���!�>��"D�z �.I��|��L��� ��«���<�~)�ꅾ�o7�����J�i�K��c�2���
��9k�Jj�Q�ks1��±�cT���d,p�_�Nq�GngF]>/�_.i���O�n�1�l+����ӽ������	33��U$�����;���6�`gB�ԳKR8�.�i�x����')�[N���l����>�����ām�
� L�O��z�Kü��@x�ͣ8E'����qo�uƵ��b�o5��W1�C6��U�U'���n��=��"q7N���3GO��N�:��l�w�m ipK��qٟI ��2/>j�p|��i�H%��Hʘ�kaflԓʭF��B��C�sS�R^\-�����g�=f��ӑ]�Ho��:4���;�D���E�S�ή/�2ߘu�ߖA�/'��&n�ݠ��H�9W�|��Z�!�Qq��q��"��R��"83�ɇI��2"���-L/9�»�^�z?F7op���l��lD~��ʶ�9%.�ۆ�����V�H-�u�hKkk¡�v��
�[7� �DVvUXf�j���v�tB��6Q�c�'B��u�yR�_	�,��Ws�Y����������
�u�3�F�� ~I/)�| �&�������k��p��t�`0�,G��B����0�/���6����!�� ]��~�%7T� �$���n�9]D�*���4��p�+�9�t�;�����o�
Lq2�Z��4�����~h���h�#$��V��i!>5���IBD$�T��W��מ ��VӐdE�p�Զ�����3��P�R���H`8�:W���3�q�-�z��,	{��0�N	���EuQ�+����k�Q���Szy}*��>K���I`�݀�ߒI�N[!]�iv�G�KF��%���認�3y-����aR��-�X�4S��x�+�,�: � 9xΒ`w�V��d"ͨ
� ����� �Mc��3�z���A��m)#[X��f���/�[p��H�~������u{�c��\���
v�{�����0<���#��Z���¡!����`+�YU�J�`�ɏpZY�\�?(�)�r2�V�^�2���&~�c"�.,���ق�`���2kr0`��o��_U�w��8+�.$���2��v?�Kb$D;V��722�Z�����]� �d�{4���+,�$̑L�3���?�±�,f�d|�H��}4�*ܽȈ��5�ƿ�8b`�:Ą0L�h`��u��V�oe��D�hܙ���_K���c��k�� �Cm�?&f�$k~$��K��C�����y��HkۻD�>&�qqo�����A�o�bo�r,<{·b��������Z1 q��g����bU\��(��.[��[S���Q���:Q�Aܒ��G���jclsa��#9:�����{��uߢ�[gς���
`y��>+�
W�u�H�q@�x�[��>l��c	�90�\@U�6O�yڈJ�G���z�:�#�"w�ښ[6�e������.x=�6PJ!���zKr�[:�-�7�z��Iw�g�pi���V�}��A�ƛ޾3�0�oE���e=Sp�ݰ�0��<�-���ܠ/�+��x=����S������I�:^r!n�d!d�?(2�bB��)�;? �
&�,�2?eiQl�S���+'ݥ�Pj�<�ot��� �&C)�� �1���,�Q�p�Y�]G�t�$� �A�|�de����z��ߗ�m��1+}�xe��[������~7Q^a��\D�7tQI����}e��l�S^BUU_�F\�Ȍ�ͭOg޹�)�#°�2Er���t!�&��j�ehb/�}��!�ك��n�Z5Z!��?�L��u#�/:dD��*���K���[�iO�-��;���rN�Ӌ'�\��]�s���=��ޟj���0!��~q���C*]oK����*�Ԏ���rd�M���r*��A�25�"J}	�D�R�+�a�Ϳ�e�G���t���Y#l's4�䫄�܁�<m�� 4��c�ľ��0�%4�86����8����A�7j���܌�3u��F�ȯ�,mb�#������5px�s-M%P&�2�L�ˌ2����7X��(���udܼ���der�p�]��X�$���*���>�ӗF�x+�a��������CZ�	8Nԥ���G�o*�Q�p���p���lŖ��ζ;�X��nG*��s�u������(u&g�	��xM1�_������'��M��j�|x�\j�:����qU#���q	c"^~�	g�G��Q�F06/K�;`��:ʠ�H��M�pKӢ�W����%
�_�5��+�
�g�@��w�>L��0�'��@�n}x�����q'��e���E�c�
郎i~5H9��GmƂ���S=W���#��rd��� 3ܩ�%�L3�n���XT!'���:��"�}{,sKa`�`[�%@���x� 	�7�>�mJqZ���H`Y"�Q�p�#��vM�O����3�n�I)���B.�r�M�Bp@��r��/~}��X�n�j�NB*���)U�=�]+0Wp�+�(�?�.�L- ��_-vj���^�!�"�]I��Q���T�?91>~(�feZ��)�˂�E��(��%Lp��3��q�*���jU�Kع�N�2[���DH��T`����G���z�S�֊�p��-%m�:�y��,Jv���1�)��(�s���n���*����;��]���9Z�������v�(�f��q�?)�� a��`��m�J�����h.��F%+P}��(G��1	�̾�Ƅ�V�WR�)��|�5�t� �l��I�{EB_7�2�yĊ��Ct�?��f��_�Va�3��݆�-�¦�:En��~un�аޢWi��Sl�����K�F�R�LW��@v�_�Bhc`P4��S}��	v�0��#/>I9�W �r�̢�=�;�j"�V�k_��;UG��o���F`�$DEq
��-�`/�P,l�se�c��N%�/tɗ�2��u�f���$�8b��Ws�Ix� `:"�Oq�r����{�gMv���ӳ�y�~��3�d^�mjEر���v9Fr�������{��Yi���O���2,ئŰV�?Q���Up*�Ӯ�����I��e�����]��K&4�k���� �D�:����&�~d8Y���	�i���c��ʃ���v�L��{<���fYWP����K+�Md����ۡ���X]�r�ɺz�}�zwc��C�o
l���&8>*�Ll�ٶz`z�^�9��&I�EV�˷�B�$!��[�a2	ч��}-��:�fo+���� <�[x�p�G����zE�o�+v4�I���@=����"�8TS	��D���,� ���_DZ�=?�PlQ���
���ҧ��qV/�L.Dk[�b�.T�B�O��!`ӟ��.Ys��3l~�H�9pu�v�-�:�~����՜�)�D�k؜J���a���|ʾq	��J�C���C�$@j��� oVQE�䎈q����m��?2��8E��e��X��~�/�d}�%�y��gn��kw�hV�}I�z]���v�a.4�"Y��H���,V>h໐7k���سI3���gp�)��}]���PhT��$�4O˭����Nt�ĕ���1S������QAӂω����,���\5�~R%ÇO=?We���8��⒧�Ҿ�r�".����	ƛ��/|BR{�%�S�I���(�q������֚f�!]o99$��������E��A֔~��\�dq�N��UA��5�?���Ô�t�#o��,8���~%�O0�ށ��`3�қ/�p�_�S�d&�9[Y���a��BDc��r"z���; eOU.^`� �5���^�VF[Ii���s�����&�k����qL-���tS`�v�}t+����@߲2}ZJ�h�����+�7�����0Ѥ��r�;{��3����B�$>��+ �n�o��FV���A�)N�!�8���WN������<t�=z�3IY4+���J}(��!�Ѷ��lu��p;�A����"����yg��s8�(�E�.�A8�/薃8F�W�3�q͌�:���`q�)di�14��se �$-�	�١��x��6�]��~O|b̪�����r�_N=�G0ۈ3|T�A��]�9<~5�A\�f�;r��6/�o�#ǈɁ	����)a�/�&���
4� �
^;{�Ev������o�_Ld@��ֵ� �x}���,���-ě]�#����%c(�2���1)	�.^p�+tr!/�Utp�3�q��+������d��L$����e9��"IcS������^�-�3�Y|��3�Wl�����d���~��<=o��4�i�[5��6��|9^��Wj7Bҕ�=�%��Jq�����Uם�#7�{�����������lQ)�X+��lf��d�<�t	Z-�77�m�_��.�ּ�(eZ�ϰ�ffi�'b^n�R�lJ����l��u(�
iR<��,��8��c*gIa�a��pg��9�\>ղ=�	NȃlL�e4eS.����f���tWy��s��o�)Ǒ�j��M^���g�� �͏Y�\(�򄵕H)��n��/�#A\#g<7J͐���B��u����g�W����۷���6@a�h��W�! ����Å����y�uN�yAN��FN\��N�M�M���,����-}��ގ�I�8�~]v^����P�whF��FP�,,��z,xvɺ�"���e���iNGP�����2�3i���RKՂi")Ƀ^�G��t��ĮD]�U��]TNXWe�>��sA��@����ſY��)��.tƧ����[��jH_�=^�ܝh���^&�i�Y6S�=u珏#]%<I�l�si:�l*,9�@@?��%�0�}���U=O1�4��!��6�q��f�{��G���EΈ�!4ܹ�A�T����.6&�֐��[��uElo�b��ٖ���d]1��t��X�t���,�>8E	�蝺[_R�~裧�������N��y���zu��_B.���L�,����'^ug�^?�'x���|NY�֣ t2"�o����aT�GE���oj)!{��4��祌^qNC�Ǌ\D�,�(Z�Y9�Q�����R���9{O�'��O��|f'�:�K�7�v?p�{M��{(�y"��� MsI۲ ��lq1�T{��V��Z�(*=�Ϋ��+dͰ�R}�f)�1�E�~��.��h�{\2��L�L�=�1�����ͨ-M];������6��q�la��y�'����X-��Z��@u��p-n#m�G}I�M��S���W��l��@��ZK݆wO��h��0�y���������Ta3�V�"������<ymSSE:��W&�՞���'+X���50Ǹ7�sȷ*�����������ciJ*S(�dϱ147͕����L7:u�A_9J�%n#�H����o���p��@�ذE�rϱ�^�6�xLfz�-N�a7�q���܁I��/��J��I�Lem.v�8\�]t=�t]u�����H;�g#$���#FKl�tox�-�����F�������ӕ:�(K �1��֖Z��H���\�z k*�$[��s�'�/,��Zz��i����7͋X�I����!5�F�P+B��UK�+�+���>ط�� �င֚ԕg��j�HWF�2:0 A����k;�h�،w=I���F�1F�T���gѽ	k�����ٰY����y?������"S�AI�<7K]l
I�L��р�~[��f!]��b�D���riz���c�� �X%����W>t1���o��]_m,�o1�ߐvz�
��Jzɢ*gL�bA$��k���ξ�-3�׋�@��⋂<XЮ�.2
U#ѫ���W~ڸP�r�:��f��^ny�\� �,��U��
e|� T����xB��OoUo ��!��>�;�X(&�W_uI���ugm�O��M�D�U[�>�ؐ����E����DB}$���]��,���n��,ʮiO��� ��T(���_�]���c1Gf6����?4���pB�9��ͥ�^���C���,��Ǟ
m��q�[��٫�B�sN�RT��f~ߘU�)@d�X�FF�K'�'�f����W7P٢����H񦮽�|o"��>�:�a�.BST|��2���FM;[A��T^&I�mDf�bx&�l{�C��DěZNt�Z.hя��g����i�� ���0�l�.+$�G��fp�͂�,	�$��R|?��ni�s!z����pD�}��w2��!�n�1-���w^�Ty�|�TKT=�|z�����lJW�.u�,btt&�w�ȑ�����8�}����y���SfnB��T]ٌ�Ԓ6I2�zE�x�Y��ܯ�8{;^�=����Uj�E��>k�0<���Ŏ+`s����(�����T%R71�Q��p��{3YĘHG�w�u��|�{Br�D�i�����o�Ig�}�$G��J��?X2'�C<���Q)S��M�J�����������:�x�n���v��䂄n��M$��S�b�-�lI*��M%/Ue�?=��k�>#s�w�;�0Or�i3}o�A$�S��X�����������K�ƶ�`�z�HQ��qi���:X�o��|��Yl��}S�5�z�5��x
�T�Ș�8*��z�:�,:��t%)~e�-d���걓h'�/�Gu��dU��^5or���E��rՔ��`C��AP�������� �4��W����f_=���uo���+�������~'_�]��HĹSH8}����n�yJ#iv ���3e`Su���Ǎ�#=r`0������˟��/��^z5t�w`,�,���HȀPHrn�����^H�B\�<�_� �yBvS�8K`&���$Nn1�,eb���L���1��\��ܲw��Ӕv���M�S��P�U��ʎ���7Կ�����]�?�(��kU��z؂�O�P����΅L�~�k��$���[�~'����b��Z2�ӗ��`����ȳ�N	��p��1�&��DF��[d C�N�oYYd���w���em���@G�t|tl�LEۜ�3J瑟1��7_Ƹ�F_4��������Tl(}��	̪����H�ɟ��וES��dQ��n��+�0eD�H��)hfV�v�h����2D�){<Ǒ�-�;(<��´���9�\fM[��+#��0p7n`q�^��8}�����[A�(�/ؚ=l�I���_.L�B���
�L+�*�GN�����tg~�ǌ�h�!3��B�<��E���\c���3�o�
i�"R��œ�¥i{c)�y�B��ɲG^�����Ș��VV�O���c��iyt:�a�$W��9m�KB�WY7|�� dR�6�
�����������)���ϗmnӌ���N��n��'��������q�W�Z�K��'����7Pk�+��P�gT�5�&�O*��d6�t��D�� ��z%�ſ�� r�~�iU+oz���!z�'��aL��^�А�ӽ���p?/����F�w�/���%�*�'�c�?uj΄㱌�2wo��|��鄣��]��Sc�xq�l�&&�@6�f�~�;���G|��ư�d��}��X�u�e���4����r�l��&/Q|[�