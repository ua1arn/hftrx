��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �����7��vc7 �pz-�0����)�|�>�Fu��a�&�sams�#���1��^�c���fFk�Ki7�#s
2zJ��9���

{�^�
\D��-�J���,v�O����e��B���?G+C�w��Z�$�+�ī#~H�f̳�H�Gtn��e8��E}Ǎ��5�Kmi����)��foޠƪ�{���N.�W�Q���'����`c#b�pj�$&g����{�|Bc�y�M�V�z�c~pÍh��X՚h�`���v4d}�zv;v�,,�z�2I�Sb����syFn�F���I�m�ۀ�F���|�h(D�t�%�Q?�!T3
I�W��<����͝p�͘C�sdP`�/&�ǚE(�WLaႣ�,q���!���@O4��
%�[LpΗ�݌[�s�G>���z��A�c��2�<�:6ֿ��,Ɏ���
�<̣eo�T���.Fo���a�����7���}	��q��g��f�B6�����{>DK��!D�4�>���^Y�CO��.�u֟��2[��f�v�����}t(�FA{��
x6^����Ody���=�d��}Pz����� �����T�.�Y�S�^��1����6
j"N\�z���݆K,����?SɋM�6S��HEu�Xݱ@g���!���V��q�.��� �(��^:��j���𿽳P䫍�����C�NI�ҁ!O5&�����	��z����=�����S@�Xl�g���,���1��@����e����H0G�(�d[�c���36���hr���7P# E7�\�%�1-c �̧P6A1� %��K>��%���~����[�U۠�^8�f��;fm_�!���.@�:V�h��X�.�m����(�׾i��Ag��ӐwQͿ��]rLM/�@�X��П��'���W�����!uO��NL�9n����158����v0u�7Z�.ۏߵ����Z笒��3:��&������EIx��K%JK�ٹ ]�~J�r-rEi�o���@��5��b�[pv�|ծ|�6��-*Rf�ʪJ�����9!lk��}��&��THA~�Br�g��/x�T��|NV�KZRux�^�W�L�7� f8�g�qbl�~ْ��Tl�&�{k ]���Њ����Gf����*�P��G���B�j;P�.����HA'�2�.%��s��ͱ�J����M)��C���:�砛J���D�	db�dU�ra�iS"�Pi3+��z�wtL\Y��)(���X;�'vW�9��d�PqE���$����bץ�䗘�|T�K��ȣl���1p���ìQ	�T�i0N��.�΋��� ��P;jʉH�Τa_$k��~��ӵ�7�9-�n!h,0��u-�A�A���l	��4���nך_ߢ8�+�%�P��J�<<����d�\��Ȗ�V�r� F]�{$�������`�u����\�@�X$��ܜ����#�*�U����c�\�N5���y�HBv�&O�&-�r����Q,��]���Sd�������6	�O�Nԁ���5�p�uۇ<��%&BL>d|�:j��{K�l���J���f�^!��[���p��L�m�����2����w��7��?.j -�V�|���"�)]�]/��	�H�9�n]�I>CS��1�p�!�K�òOL�e�c�7}�@��������ou������,�S1��A���}A~�1f>�]�X��T\�g0"-i��Fq��\��=�R���j��H"#=���O�Wܡ��k�ݏ�����h��6C�����U�Axx�"R&Ч�֐g߷Z��Q:����^m>����T!�C��"����խɒ�O���z�ai�&��W�1��L�� &e$)������.)-� |��oe�K_� �#��[)E��L!g��/4\�3-|(�T�存��+#x�QB�� ��F�!��!�Z�&��8��{?|�H��;�b)ځQ�"��=1Og�j��ݱQZУ�\[5�x���� 0��� �L��Ġ���[��ަ
�q�Q�*UR"L�mE���s�$��l۩6)��Ch�#�J�}&�Ǚ���u��MT�R;y�d���}���[57S�,��$:���`�W�S���_K.Q���Qx���'�B�;��Js_��Q���f�Lj��H�g<A�^-`��t
֭�ߌ�MDFY�r1����@7(��)���PFc�Ef���[����`�i�yN�MG�'bVɜ���K�A\�k��.{���'��҉DF�9�n�jg�����E:t�tX�9�q`��װ��-do5�/Z	�X�S��~���4��)փ��+���<��r�z7�EWwP̪�闍��Y17�q�ܞ��̍6���������Q{�U���`�ܫu���.��|PX#Ady''�!����i�8���>��Q�o]�ѩ��x?$߶H���j��/Xޘ��7���N:j;a��!ײ��&�}��f�z����-��w:��d��Ja���͸j�iV۵R���{BKp�a�c�l��],F�&ur��R��������8��Γ]��1�/bF�OIH�   �/�g��~��î�6ޡ⃻�}SV͝Ǯ��*��v)��Y=�(����׼̡��Q9���b��-��ɐ�ϔ>B�a�`�㛶�^%Pnbω�d�n|Η:vaIԲ��њs�M,^��4�p�FfR��!����������u��q�Jsd;�$7���?�W�)P�SO�'<|q��m��kP	�����P�ImA��Ո�:�*+�,aA�{k�����;
�%\�%��[Rnɱ�&����S��丠"�R��]�lr��	�h�$r7_u�g15��3��7a���Hh���;O�2� 9���!n|��E6����������݋��V߀�B� �ғ�+�A/Y�Q|������4�9v����ޙ�E��Ҧ<�+k)߉�����7'r��W��l�.MIѢ��)[�m\zQ{�%��ãn�ZJ�.�d���e�
�{J�@�P��m�	Z%�u,�Z�'Hub�����[��������8���v@5��Խ?��~$
`���o%]�6Q'��Њ�7�-˭�dt=g�!5�����A�ݗ[����hԪZ-��4��ӿ�D!ߪ�+->k�3����J���+2� �g�����d�4>��(��,a?��3��{�g�������,%�W���/B�5V��j�}�X&��1�?̑�ǌ��*ߋ���"q�[��U�v�\���Mt"��d�sT(��A��%���XJ���jo����8�Ǿ�B���ɔ�1�&Bh�,��N�����ޏ���3�!,�	�ˬ"�3���ʬdu{������["�w�]�߬�i'0����p��TY/iR��<��9��¦��F R���w<���S���V@� �4���D-��>�4�}H� ),IRgUF��k�	��T���-�qx��CA�<�=����6Y]����`|�
TI2�
��x���i�q_�_��W�5o��E���d�Y][��z�/|K(Ij����y0�*Ӣ�
�B���U
��y����O�TK|�U���+F�[���Չg��M�v�7��&I��/�t��H�t���|��:�"W������%tl���P\Ь����I��hqCf�L��ũ�
�ܮ����S���d�4��v�G�-�͓�e�k+CӐ����w�����g����Zn��?ꃇ˾�4kz����9K|&����w�"�kS�|�1yNY&�Y<�����.� ��ݝM#�"�J �2i�ZB�P��t馉�(C���<��mC�}T�9}��SB�*ZY�}���V<�N�̤��˿�Aޙ� �Et����.N����H�i��EwI���MJ(0+����kk���U���\ZDS)jh>6����p��giO$����$�+a�̻Wa"�"6$YIW���)@h����$�f+�d��>��͞�D�������n�r�w;0����u� ��0:�u�2H����-ʬ��I��J��up��}�xw�K��h3?��Pϗ��i���\�fy��!��Y�����#{:B	y���v��$�����0z�T+�4�}[����_L��`�����
c�k�� ������o�!�Ơv.N�'� �A�!�i���*���/Y������ȍ�.�`��(K��D����!k�^8v�N8�L*�5;O��TM
��wx`9���v�F힉cjPx���K�qw݊$��#ۉ�G�����lpHs����ª����8���C��]��
��w�Oڈ����$�2���ن |�ٵl���b�.ZȜٿi�vƬk��j+��I�e�3����3����-��6RU��K^��G�oJ��OA��/�%A2�dqY�7���*�+�9�p���%��Kcw^
.ãZ�8�iq�tؤߪ��뼟�9d�����	�\V�l�J8a$�E�;�V@�A{.R����-� �z&s��p0؋i��*K
O;k�I��~��L:�S����j:�W�k@��Қ�,�� 8�>��E���)v����H��`��pͱB���5(j,6c�2 /3�~^�Z~IϜ(R�K��玍JKdB�;��:1���A�Y7�b�����\+�<K�]�wW%T�7�ph�=�ϓXS�m?�D��SϮ�����*rMQ���kԲ���y/_�	����v)��k���#����G����ŧ?�ɜ�TO5ЉM�yL:��w����g\+��g�U>�����t�8S��#e3��� ��6��n�#͖x������y���@�R��5���L}�u�ɱ���"����׭���]�g��/�>t��w�2��L'�4 ��r"�^~�[��o�t���oRkFQ��J��i�_ t1@�B��r��>�̀��I}y�� �oafȾ!��h��t�Մ����������U>�i��K�fC����ﺑ�A���Wg_N����w��H�*��C�x
 ���W�n�"�ۛ�5��%	����4�Bm���D�À@.�2�����Qٸř�Yn���p]�s]�Fx�FaB���c�4qQ�'�[��P�5�bg󤡟�Kc������4��i&�� ���h��MJ��KW���0��?TdU��ǐ��$�	�� �&K�Tu���j��)g����hi{��֨ƛ1n�I���$�X�J��V{	."~G�5Æ��Fw���z&�'tA��"�c���w�&k�:_��u62�z11�g��,����ZL����,M�����J�;��r�.�!=�G�l�[2��V��fTj^�LV��	gv��k0���<Ex�R:�`�U��9��7s��d�ss�O�%�A��U���dL�����+.?"��F{�lA+����za�
�9��^Rǌ![���؟3:���<M<%buH%��U��/.T����JhA����X_+*}�gx�R0a��'�6��M��Ҝ�X�ضEʼ�H���l>�#ՕG9�4���N�G��G�뿚P����>�W �c��p�оd�q��Y�-��,��G����k�N/I��B_}�:M� hK�2��$)��^�m�j��>`(�p��@:����e��?�QG8��=(I�����f�P��+4e�D���8��xf�\1�fcO��>[9o�9�����#^�C�O�Q��enw���Ar�<��������y{	ZM��s��)�3���B2*��� �*�a���Ʌ����*��q�#� p�T�Y�x�MHq����>.]�7I~�_�9?��R�7���"��M��%�!5zQB��c����ī�~��?���������s���<Ի��Vz�'N�E�)|���;����#����9���|g�y�p?P���ly)��G�@>w��`4�!,�!��m�Cd�L�����c��/��9����������g���>�Gʆ�	#��]�[�t6Ò�'3�<����~!������>ㇴ�5��d�>�ėF�t����x��	��{�J*�s{KB���2�|�x��王�F��D/o�Bf��%n?��7��ڽbȮg\�_~������ax�Q�d� c4�A����IɭG��L}������!��W���}d�;X��}aZ➹��	�՜���{�H���ϱj�X�"P�4��q/ϟ1��rF�(E
����G�5�5�G��Q��vw�i�rbNh���3�U�!�uk��@I�,���@���Z��Rx�U�DCW`����0x� e����� �g)��o^�zƉ����܄�;N�r�|�J?��I�����$k��:4�k�q��JKK�r��������y��5c����_��u�DRU�K�6�t�~����h�h�Y�S�#1�~�Do�b�Z~k��Jj-O�e9�L���Ͽ f��:��
\���ȑ�-�*d�X���ͭȞ8Y<7�V��]��-j7֪�a����NL�A�}6C���`Shoa9�K�WFMm��kȁ%��vg#�� ��ˤ�I�XQsR������b˲��q��`�}��9��,[?��9�N+ $��9	,��<T�<���,[����Rh�a���@ ��"�+��,���J��7��i ik�����)Oh�����&_�:���t���u��)~����5�5���伛��ьo�RFҼ_���
�K���/]a4*t�ڹ!� �.Tu`�ڹ\��sOV�bEZQ���/p�F �q7y�
��3CJ��; K`�B�C�2ɭ��9Ml�����z|��k-_�O;�9x�t�����4�3���B.�����r��C�Pc���sN���Y��C W�s�U�`3��	95��AX�F뗭I'}u�?6B�vi�2�����呍\y��W Y�a,]-���>=�[c���&-@9�	�()�d��n��n��P�������?�l�Z��b=Q�pV������;$�
u]z4�����l��h���8s@{i�Żf��qU�;�*nZ7#D�6�ܠe��җ{��e��қ!�����1�h�n�l�G��I�I	�ɬK�͂P��]�
̧u﫯��/�:�RO U�<1 �\>�ߨrQ����먯5/�68G·�e�v�:ɋ�2��P�|�p���+��G���������[m#��k����1���ȴ��}A1�����>�Ұ�-1�	����d���nٜFQ���+�����ϔR(�l`7AĔ�|�A�9Vɒ�ϲ�A�C�\��w+`�=k�;lrH�&�\Y�B$�����+_VNUo��d�hu�d���
Ls�	ɁFku�����x!��d�����{xɵ+��p��$%hW��� F�$��&Z�\����S��-1�O�~�,�����䅓�̞�X��Q���-<E�赪s�7*<�iy� �l?�Y��8U�t�^��(@|�#p���u�%�ɹH�%N����E��ȥ����(iuo2���SZB��ޟ6���v�y�Up\���/�:늵	�(ȼ�t{E�X4�����F-ZZ9�%�a9�o8�/9�K&"ҫϯ��=�'��o��M$uĜe0�8��� ��O�rF��/Vs�=pJK�Q�3m)����_�������w���ٷ�t�r(�x":�_��Ƴkj�MK�I�vRp%׭��45!�x��1��C|���$W�w6$�tD%�HykI����u��$Z[�Ub��φ[����MR!��~JNU��֏R7�Л��?2N���� ��(Ѳ�	���IT9H�$�sc���.�5T���5:rF,tYK���g��?3;���|mh�q�/��.;5��_���A(L`����&�!Ϙ�fbR�*���Q����_������B#1��"�#�De�S]F�*R���+*�ֈ���|%����s�}�`CQ.�YRS^$i,�*������<�����E�Ҁƽ*ʮ�$^��Ku���A����hj-7m}�I����΍�����N�r"c[Z��:�Y���A�\o6��|���DB�~\��g���t.UԴz�R��~�t�LuKn�^�g!��/�?"o����I4DZH�Ib�o�:y���I�4�#x�\���,�6��GP��,������2{�$ajШ�P�N/!Z7���yÓa�f�VΫ�0����)�uw��$�[}�x�]Z���-�U��p3}��$j��uI�8�J�d�J� m%gq�Ԣ��G��8d���~���n�U��9ÑXN.ʂg�Y~��2�#jݴ�����<Z�$�8�&���\�iC�(��*��V��)�3�??/M�g;{�w[I�NEu���1u��7�Lw!��d�Ԩ���$9g��L7����C���hl/3�T8w�������|+}H�uF+@�O�"̥�]e��I��=��]�O�p�h7a�z�����(��z��@�g���}D�C7r��-���&H�c�:Y����z�9�N�?b����A�<�L���L����^Q��!7$q��������&�#�c��M�`�uN�ǈz��Ν��`�r��9"�MuU6��%���sfOz��7��]�u���7�8�@Â9}����;��<t�k�2k���W�@1LP@�v9��A6+A(��Ց��;�g�������l&�|[\��$JA����,7��_���x�=�~�PFQ��i���I��oUc���"S���(��j�h�&/���d3����<m��Vɝ��CT��!���D��k���K�+����	�
 ��71�����^Y�sh؛��DU��b�*j��&$����,���R/�\ۀ���酡���K��u�s�"ЀЃv_��xn��S��S]@O ̈�M�-���zb���X�s�s�W��!���e>��Q�}��J8���`���/�rN�{�s��b����uvE��E��Z�;��+���\~�u'��op�GI3�?�|� 3ȳ�G[��uYp�킜e�2҄E�X(�E=�>u���� �q�l>w�Zɴ/߭��Hqutt�--S��F��Ps��8	��&ؗ����N���V�3�@�yT�)(��#�F�Ď���r��E�W+Q�4�D�q�9�")�i��ы�N�;���|�O��S���D	:#;-M���ARt t�J2�E�i���HK���L"*���:� ���FX��⿚��eR��W��>� p�z/�N,�H�7����x,`�&�+6�܉٫�NkÛW�ҙJ��5BX85����7
-͆��A�tZQht�xi��~�i�����b��}���C��4�T���utscu�-�{�VSV���qI��݊��&"��-����\�G��)��������<]Pvgp�g�P
@�%׆��<L��� Y��;�lTɡ�GpH1�q"��u��y3�{��V�q�<w�kٴ���V�au��Mm�H�ˇ�a��8�� ‾o$W�ٸ?�z�HN
���mY���|��|
ȴ%����"��z<������퇘���LY��P{"���m���}�����֓��D` �Ѱ���.༅Yt+O��j���E�_���8D_���:��k�J�n�j[9�j�e�VA��u>4u!d�� ��Я���X�^2�Ӊ V"H�W�b�	J���'�f������'W�\�J�´j��{�D�c�L��&0ˇ�pvZJ�_���P�l)Ӏ��anx�>)�>[h�]�i��1�7]C�z�5/��h�V(K�>D�C<'��3����K�(�$��2"�7��E1����\a��3.�[Ve�6���_Hg������On�u��/~��9�R�����m+� U|����MƜ�qg��@�O���ы�N���U�1�z8OȆ����:̒N�`9I������.2����J�ǡЏ��B�cȕ
E��<�-�q��Z<L3ܛ.[��"^�?|�E��L�u�Q�ݛ��z�*6Q�鳯B�$Κ�ԏDu<�?�xz
����N�dl��D�ٹze;��5���=����*G�ل��|�?���Ek7��d_�b��d�s]�Py�7%�7��c������O ���]Epɮ�J1hl����K�1ݩ=g�i����v�����R��/�n�'T�	�I��/D��

�p�����>�b,Nޝ�ssC��T�$�!�u�WX%�ʩm9�+��m*�L�W�Y�&Cc؎s�߶���Y��J�(��j���}�O�a���1�#��B3R����O�G>����+�{�v<��P�:�'+���"�t�X�Y��o��� �f�d�h�e��^��%��>L�)�Ӝ�f����G��7bӣT.#|J)?�7,���'�����]ȫc�/��,��?�*="�<,qQ���g�T�w�!yy��h�$�GX�[�(k_Q2K�E-"p` ����Uņ��vBA-X�m6��4�0ͧ�3;`-�Q.۾#�;=3�Ń�ڋF�l���ՎF� �!l~*&�t�KS?��.��*dy���C3o�'a��^d����PI8,���T�1�p��j�H�b�������J��aYx�D�^ժ����{2�vɭhހ�?|CA�q)er�_JBQ��ݥU/���f����K���"�Е���p��ŵE���lӂ�ŷ��Q�El��}O������UA`�bi,�r{�`v"����Rs�Hr��૟ܠҳ\�b� j&u86Qg�|��q8'�H,g��.x�Y�Kf! �����p���t����'� `�=D=A��ܢ#Q���.UZ�!-�s��+�!��+�w��Ъ��vU��W�1ƌZ�Ҳ�A���,D.�c���c��S��d��;��ԟ�]����j1�*/�� x�N�������R?v�	����I�Z���F|��%��:��87YU�`����كf#&h���npX�1'���c����iXZ\�EWr%/�_c'���<��2D,�U�x�8Mf)�L�'������%�DS��!۲׽E!���c��B�+�^_E��F'��x�*�d�cF��=ԯRV�2�Z�G�(���e�Ʊ���S��r�/�U���o��u���߲�O3�R0U�|�H�+���[U�Ba<��3��ֶ,�r��h���=x�5~�"0�ہ�X-��H������E�j^��~����Yt�-�3�`�%#���Zo�B䳊�oIV'��H1�vl�$�sX1���m�^�������k�C<rq���!��ծt1X@�eU�5�8�Z�(�-��&�<�����7���T`�VT�n�Е��&vs��⺢ۖZ�"�u���D5Q1;R�l�2D,Ѐ�c�`�ӪP�Ǆ�n��!ǒ�0Va�=me �=�IR��md`�.��M�4���5���Ἱ{�+XR�1Z��(tc�Qbr��l_7I�J�8��-��V1T+$�
Y|��%�+|4��y;�F	�M�	BG�^_a�)o����;�������P������?��_\�OQ���oP0�5�Y�Yv�.y6܋��,�~n���^��������:9�6!+$%"|�]F9d����[��hٮu90ss�l�w؈K�	4®h���= .��/t�a���vL�b���;f>�������h�T1���:����J��s���Tչ8B�7�8�d��㻍;�N��D��H��ş<��y��;h
�^�iQ-�����=�m��c���F��5�Ω�Y��n��l�!#���t~Ki:�-ڈ��b�7/�����^�'�?]��-_yp���ES�UN�k#�����Os���5�3�@����;��θ"����nF��K�>']i��\9��n���z��haC�S�Q5�΅�.	���e�x�^�H֓�8���>����7^:~�c��1�O�R�]n�����g��&1�/�o�:��=-2�QC�W5���=H��vE��-җg�&�f���4�9Fe=�m~T3��b���� ֏�FL�)��P&�s�H	�F�>6}�j�c��ND��7��=�|���hP�Z���T��>��[�>~�)���_;��<��pה�C���:��[�O��
ܠ�ǧ�`�`�?�}�]-��?���դ �l�m�y���#�idH�|�d�Y���LP/�;�����Z&��ll���?v*��<<�<|���#�y�m�B}BOϽ+/̙wK�1� X�g�n`ڞ�E�I�(����2�ni�7�h�s�
xI`3�����("R'���ֽ�`?�`��o��KOƤ���綴��I�\A��Ϝ͚~z�݃sA���`����/���	�C�v��:9N���� �9�<0��r0�*�� �I^�EIܡ:wf:�Ph
B�[��&�w�}��h��Y~4��lsJ gv��U�/��Kˑ�e����P0sZ�Wk{7�T}�]I,��iN�9F��<�]��q�s�fC�|��ER��vO�(����_j�Ȅ���Z�����yY��{vbUR���N��ڍ�Q�Rq��Cs<|�~�-���sm�k%�Җ�Q��,4�酁�|���כo�bD�S�cv!��n�S�jM�|�Q$��P7��.�6B�҉w�Q2O���j쫬·�Q��S$(��b9�~t�q@���z4�*4;��)���M�t��]�$1u5�@�µ8K� 0#΂z��z��NBВ�&'^ -�Zj_�>YA���e�GS�)�`V"�$���?M�xn���:�7�����\/��JD����X";OU@3����E9���$�B��XA*�M�����!�I -���Ţ������$��S����s��7�:y�}I���QC��
h7X!�݋���
�G���3K�f5i�pn�V5#��;!)��ވ�r��;���&셛 TY�!��dы ��.����+pi�6��/DD��h������D�U��q?/A�먘�'��	�~�R�	~�� �G����g/����i�0*�QX�D����r��©��qqyj��_a+;kD�����ø9D'hi�u����g =�����j���}!�}sa���-:�� ͅM
��]�7fg)O�\���ȎS���K6���7�^�/�`֔��')��dG�Szߛ�?�3�m4�����8�y�}�Q�c}�M��[0�Y ^v�x���Ȁ甩O��
���2\�q=<<��3j7k~]�����X�$�Io0d�Y<a:ˤ�C��ei�Z{,@nB�,P�ʔ��DG'[ER�np��A��#��\� �G2�,�O,�ԏl�h`��&&���(�EA�S�-��5�^'E_rrx��iG����p���lսV^ �հʴ��e^{�?3좙_A+C�!�ʸVy�<���m�%8�&�x+�W�\��u��$u��FԏO{��4!�|��?X�׻ݠ?Xz	�n�H#>#U0��s(,�>�b�Z�Ȑ٭����{ 
�j�D`�=I��c��A�q��m�X��n�]�aa�Ԩψ��S3�@�����{D\���l���j�B����H-fyQ�3bġ�=ۈí�����k>�±\Q'N����2�r$0�~��D���y6'��<��a��O[8���M�+�������-N���
����m�4L��kw���0*Uԕ9#�7,H�W}�YP�W��a'����EѰ�XZz*a����`�_�ǒx+F\�GFAԌv�����)4 _���쨨7f R�"7�,Ph�`�U��k�Mo0�a�k`�(�1t}��`1��u�H�^T�?����5w��a�_Y�2�S����ԏ�������t/t�U\���JKٵG��0���Vg9GFY�=�k��BѦx�W	z	J��T�M���\��I�Kմ�`�(��Z5��7m7��3=���P����&�'�E^��w�k�������(8����ˑW��&EޚO���]��T����J�>��:�BM"tӓs��N!��+'9H�ϓ���s%8�a]�hB+��9�h�iO��Vp��^60Y��AX�xf9ݖH�$�-j�́��]�ȘxU``M�d5�T��*�����.�U�vsO�h߱��F�+2t�coSB�M]���*�3��}��Q²��&�7�0K���d�k}zP[ۭ��O����y��{� z�F������&j51���M���o�+z��A.�q�CD��0���LZ��j'{޲��h�,���4�G�CoO���.��t5��z|r]��0�8�s����9Z��n� `�p�QDO�V�#T�yX��w�N�ϲI�q W�5�>]!gH4�8[�xM��мg���h��lέF��J���N[�1�ȗZG~a��һe�	��;��*^i7ݒ��g��<���1����X��݌배���İk��Wn�g�OPM���jk$��o�?�k�A�]\Vஜc�@/v�i|U�s�G�v��n�����?/�A��<�t��0>�T�6HU���m�!>���n�{I�1���6W��6נ:tdo� ܈���1��D�@�����
=�=8�t4�;�4�`z��c���D�ë���֙��~:�v)"!�����k�M-<L�G ���7h�M�G��b��^��r��uK��jQ��3%*3�UUAI�KM�(Yz5��?�o��L �9��xh�P�UDa]�O�����C������Dj�ю3�JT��d98�����Lhe�9r~�{hu2�G�k035��NnE}�3(#뒸����Z�5Tk	���{آ«�c��K�Ŋ�F�����p�������}w����U{��!��ʂU� �vm��e��ӻ~ 9N�sx��.����4���1)��#Q'�G�#��������
cV�r�U:οv�῿�HX)̏tP�!g�	�r���$�(}���YYD4M��uks����8�z�sF%��Wj�>`�#�Oޓ�gUP�9�x}��+�$5_ƣ�#��k�&�����`%� �N���ړ����'+̺ E*��O4�֍W�5�C�E��q;(��,�H��;'����<L�%`��Bd&�q���]%�"{yz�j����pP(;��-���F@���gO"Q��6��8P����)�t"�n�MU�=(β�J�i�����o���l���N*�5��/>��;k�����ջ�������-���+�?��׫�dnT\�UA��uCh݄����Z�鯯���X%�Kd��ټ���=xĳ�?�9�H�T<����5� �����i�,=n�)�������	(e��X(V�C��`«��2%ͶM���C�Pp��7�"�Z3��!���/7��L���+�^��&�V_�H���_��:�Q:��������� �DԜ���%/=���Z��l����n�d+W����6��x��K��4|{ǁqh���6b����xmS�ܲ4�J�b@�Ĉm�q����Ɵ56V �AI�&���U�|�� ��hꃨ�U0b��7�]�{V羍��3Gܸ$hN�B�i�j��G���)�Fޕπd�����w�[0`���ӈjG��|Pys�+|0	��;��튇^�BT,�8Ļ�	P9�̬j�w��EŖ�B�ح
�ĥ]1T����� �Z�x�Z��*���Ү���Db�\��@���	��O��j���L�����ʜ��#�B >��37��E���7sxx��R�G����v�����g�7:��ͥ��۔�1-A��_���RE�f!�/c���CTaM��We��?#l�Tb�F�ZO$���ʚ�j��s�uԗ�<<Æ�::��;����l���E6�5�=�a�./�}��71�[TI�n:`b��a������^&|��m!`��`��L�@lV����g�n'�A��|��U��t���	�������V�Mā!n��Ƹ�!��ߨ��:0xhe���S ?�yp_>�y��e�g~aHaTD"	��P3�h��U%����^��q��0���JT��h>P��ٙ�K���
�M������><$|ym��O���*�\���C����O���|E��8�߿A�]�O�9�P�@�D{顖�y/Iq���o���אk>���9ߕ��|�@�;QEt81��ti��Tc��܁M���H�wݐ.+�.�_�ăY�Y���<�$�D{~rg҄o(:x�����O�H��=�O�6}y1�*��� }�;#�1���"d`Q���ɚm�����#�KD2�_L��:7u���k���;k���jT���dg�����%�X����y�u,��qq�v�-�j�hNaPC'��`��,�1ܠ�P1ׁ��Ƿ���	��?��������S�#`{[�����3�]|m��*K�\�E @�(�*�M6̛�l��NF�;��R��5�#/k}9�t��ڍuT��Nl}�o3)6�I��E8�F�"�l	n�>g;�}8�A�[�LI��i�����7�c=p`
��_�g�D24�=��)s�Sl!B���+��B#Г�L���}����~/�F[T�"���2)��⑘��z+��C�^�^m�'��;�^'�4+�]Fhhd�P�"|���!{�El7:�kw+`�"�C��\_q��SU��@ř��UO�����K�
�������@U�$���.�jH{T�Τ��� IZ@�+��h�-Dwz���9
�$-swg���*Ԩ'HJ;+��
�F�qZU��|���/R����֜皦���\~أC�:��i|d}�{~i�~��W.1(yE�װ�Kq�`u2���9թ�mK�~��s��>�������8�3���
���%�f����<%8yGׇ{C�4#	��I���ԍʬ��f�F�J�u+��
�X�K�hX9sQ�B�K�9�ZW:4u���ݡ���0B4:�׷�ʬy)��ډ����A�4j����jD#��A��l�����ׂVG)�� ��]��Z�Hs�Q��}용ޜ�#�D�"�5�5蟝�z��68>z��㞼�麚lc���5Tag9-��D�����i��V\�;�P�z�b�'>FY��0)�ɜ�e��*��Q���N��4�]E6;��쮆F��Sϴ��n�u��Yǋ����f���? ���H\;��M���0%�)�p	�'*������A`��,>�1@R���
Q�7�c	q]]ﵱ8�v~#�Zob�P]��(�\>op�F(����p����j�T���S�0�\�JY�
�2�5k�4�\l"�Z>�}��9 �P���7K��;#v�>��BO~���_��`�+��G���%Һ��V��CsO��mn�,�֚����*&��q[B�̦��n�����k�,aс?/C�|���Z����?JJ�v�~CH��1���U��\b�ҥ���"Ȳ�s�1;Jε�4�����#��P?Sr�7u9�jS�N���*�(�5F�޼T�K�`8��ȼ|R-5�3�iso�]"_����C�.%���IR�*^�����x��pD[T�]��}6 �c�s��B�j�s�P���0��"z66(+?���'��&��x!���o��1��a�-�"S��"��T�F�"��;�F&���1����;���(�d������rc��Rhb�`�EsIf��Ӿ�l/�5���[A�lh�c3���S+D���^����(��$6H����
�8���ntY0$ ����M�ߛ����FC=ȿ/��}��r6HǶa��Z��$�|WI廐FӲK�����:�^U��D0��Q��B!�,���y^'5�d]k\��d��^o�I��������A%�=^�_�E;�g���a1Р�	]4;i�wH�C��gD��%$�].H�ԩ"͠��WF`�	'.l0���H)�Ų/Ⱥ�P�oOԑ�4�|[� C6N�w\�>�����ps	P
�I){�&�@���ܽ[w�S�.Q�>��3Q~�_�"CY+>����q���g���v��CL�.�Ao��w��%��>�[�P���<[��(��:v	vP.�����,�!O���T<40�o�ǟB׀8�5��k�d���m�R�>WCC�H0C�VA���F�^���_bt�Ab��Pˣ��>����Z����Q|�߯���
���2�/�������c�"��=�UB���ԯj� W)������r�3�ր��'7̤ed� �,i�����.6sԮ��e��:�f�ULP�U�-���-4�������*�2�3;�QN)�x�r����"����)GBW��J�v�ֱ3B���V�"��?%ҚhtE���^�YI�$.�Gi;�(<>i.�϶��~�@,F��|~��cy����a���^s��Na�����Rj�o�k,� �+W��e�����s��]K��8�(�ٳ��c&�@���T����tv�����DpZ#�������H�T����R8ʏG-#�
�T~����%�_�7y����ҹ5��7�6]��_��]���g���fo�>�z���h¬�fُ6P��ϧ ����џ��5���P���4��1�
��d�+�[��l(gEKM/�w��~�ɒ=X�*$j ��>�t\��3z�`�ҀQ�j���S ̉N�����p..�r�h�Tf4��|X�  ��<��r_��[��(T�A�l#j)�T�TO���ߒ���j���Զ>�'�if1n�%G��A�]n?�E@�%�y�e����*V���+�.h����q0S)�ل������`ء�3.��s-�,`�(Ɩ�9I
�����<"�Yъ��E�I�"]�@����Z&(�*�FY|4w��w�]�6���sCS��s��A�$=�T� J�b�`��f��}��6��L���4vt����s�H�.�M&�H}��7uVk�!�a�a�-,=�f|~Xmu����5�y�	n��_��h�C�_����ܗ��y�M�V�)љK�:�2X<VՌ?(�1D�1 �:���f���˸��+>VA%K�MR�_F&�c�U�w�h���ݙ���oGt7�t\l�G�h��74����M�#cu�G�x��~����`�]��޷�wX�G�*��-��7���WbA�/���H�Մ[*�m�햜���d-/"�kA�$}�_.vu��`��%�-�['f�Z����~�{���������z�^��������e�<��6-/��Zh��u�8	��ZNII���<�/W��|/�5e�L�8$�u����B�������f>�%�[ Uy*�^�-�dDꚩ�33J�3S�!�D�C��h�;�bg_��_W):#qCY�yp/Y�U�F ����
�t�V��'���.���y�;j�B]�$�$S�G�':}n�u^0����Tv9�|�����{�n�'@��q�����rK�[z��tsdb�^D�><�Q'5&0�j`�<�M^芴�ر�!=Z�ڷ�lO�F�%a��}�zc(��K�֜�q@���<A@��ܷ}Ol��g��ЀI��W��%�������8��T�gq��V�@�6�B:?{����g�`�o�\�
o�E2�bF��1(���g��W<g�ÄZXHՁw��DN��mM(�����S�)y�7b78�Ź�]��������?f��V,ei��O�~`5�ؼR�0��&�?*��T_?��!S+���2
�����:!�m�k�Z3)=��_,�h��9��&m�y��h�_�Ud�?
�&�a?s��1B�w�dm��H��2�^�x8�uI:y<�~B�%@��°{�;�!�����q�i�FC��2��в����U����-��G>��2�T������Y��)&Jډ7.c���숍�gz���~G9�J��a]���Q��W3�I��X�S�L�I��X42J%�@  �묙#K�S�˅4�zö�@�w�]Q�n�9n�}*�Ħ�?���ձ��2��n}���l�ŝB�R��mѨp�Gc�o�k�� A7wr��Ւ� z\k�B �(y��2�5��^�I���.d�~�;5&v��nQ-4��=u�m�����e�:�߼۱��q&���.�68:�P��n_��Ma+�6�	���F*��u4���2�3���ce$M�[A��8�Ǉ�TN��a��?s�r�U���e�PIo��Æ�'�����t����X�;ů��*��9%�$�+�Y!��-d�g_� d��.%�%l2li�t�*� ��^,���"k�����ih"[�o�'x���0 _��x8�q��Z�=�x�7���3��/������ʡT�4��b����S��IG�r��c5�[�����u�>��#B�2>l�#)�L+}��Zuj�J5ՀG�,r����&T,�L�u0�#
o�`k+'E���,h	��B�ǿ�sl�.�y�����~���Q/xFRߥ���'gPc�[�+��e�~Fh�Q�&R"�0]��*0��e��E��G�}��+	�T�L2�j)�ל��� ��E�B��9b�m�-�C�F���P6N�e.��
�`�q;,y���!��|�R)�ǛW���kt�����C�A�(2d�ÿ�(��Q_��x��I|LA]b�G�2��Lf��	I��!�r|ۺ���*��g��@�ab��1��Ȼ�쪐z;���-z�4��yv~��C����\���O�g��W<I��M�1-l��@ӚQ�,CC�+`� t[�k�K�<�ㄮ��w������V�ƣ���t�6��_!���hB��3�<u<���c1��6��r�ڞ�DW���E��JӿP�7V[b�uU|+zP��h�a<t����9p�B�N���#翙�O 󾰹�+�}��a����?y�3�� /��<l�^��5u�G�q_�G4�����BrH�՛��,Y�����f8�{�Sd��ɚ�jC���s���)��>����#�тc�4�rMyh�Q��cf�,-`���av�h�1�?1� ���-�� R;����e6�E�]���J"i�b��f�\�3sGZ��~�a��Ce�G�ڽ��vV��q��r��b�!c���W}�UU%�u��yP�E���ZȈ�ò��ߡ��\;>���O��?nrʁ���tm�N�ȅ�a�K�+e��t��ݜ��x3�ս,�md��ˢ��+��HL#k���Wl��E��|H*�6)_I�S��j~���cM$ю�:g�'ٮ0�}�柆?��q�'d�E��b����^�@犡c�1"����nBx�ݣ��㎊)�_�%�i/=�#������E�Zlj���h�:�Cf����*�����zp�:XQW��
�ugCF�'a�g��M���
��;�����NfU��T�I�}�<�/� ����ǿ�F�! ��u)qb�s3�u#�ÒYH]Q�؇!T}���t*��U�%Vn��3�O){�����@E^7�b�X�JҰ�QH�z̿e�=�k"�Ck�qS�DB�DH��3i�9d��q:�nBʃ�dV�z�|iJ�D�{Z)$aE�P��<��ॏAT��p�0������p4Ȟ��<��+�S��6s���+�+�*���R�+��sNÜ<�0�����J�NS��_D���obo���c÷�0�2�<�&�� *uN��M�Kz�2����P��A��%�۸M;9T�it%��:?��~�.�<e�kv����C�Z�����BSM�:p����}��e��"&):���H�H�o��Bk�m�R��vP$@��^�_����e:��U�oq���=�������)Kg4gEM�H.������$Dک�abk-Y�:0Ts�����^�7��q[��(��o �JjJ)�gu�gM=�*m��g��cݽ׷2�&7��a4v%0-N��@�������gޥi��p�s\��1N@��-�B�7섔���� ~���d6�7���J^Y���BO�n.���%l7�ۗ�y��_z�e��C��P�f�m��
�P��JT`�����,5\�-!�hr���+"�0���`�Zp��[�t��#C��pu���a���owEy�|.�lZP0��]2ݡ���.���ĔL�C��֒muId��x֕}T �&���K�WXQo��t�Tr���|���-���e��æ���p<���k��|��"׽p뚤$"�M��$Q� ��K�X+W^�u�l�	U�o��}AopZ��/*/���M񻌆�D.�����9X"�1T�Ą6�ĹQ��D}��'qD*~ϼ�J0z)/��u�����<����H�ELM���Ψ>��!�-?�"��	ːhS�������Y�/�Z*�-(F3'"�qx2Y:s�N7g����R�WJ�^��ǹ+|�Gv]��{>7Q�����+Tc��v