��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+"�:%V_��	�Ξ�܉�����_̯��֛%�����A�Y��Y]b������ju��e�c"Vo�32a�_�$�X<#��7r�C��ڳ���Zm�^�@��!���x���E��&2R��n���{~[����'�Jտ�P-�"��y�v�L<,FTJ4��8��ŗH��]K�Y��q��+B���;K����TI����B�̤
�S�!�QW��(x���IVYZY��'���/� �;�ݑW�_�'����΄
+!�����yÆq��1��.^ݷ�:����΁�RZ�*gP��E��@��N�M_����=��B�m�h�b��Ē�I�W�b!��+�VU�YV�� /=���/�p����洆W��n�Z#�Al�^�L_�=nv̆������$ZWP6��H��6Tn��k�5<۪jk�hUf�mu��g�V��[FM���ikZ!?��̪=���n�$�?;b�k%��i(��?$f@o�/�\�H���5r��}r����/7�ê��.4��r�2ES�R����7���vw��P~>U�C���L}dy�ToG����Z�I���W3g�qcs��$���А9��-Yyp�7�ċ-������\��@X�XD����p��ON��D�T���[��ř����.�<vI������}t��`���q�}1�%l4ê�[l���U�"V9�y��'ac2M5�c��v���HA���6���.6n�X�$�dHg EHlH��6�j�ݯ�
��?m���לi����\ru�U6+�TM>M�@��we��D�;\z�]:Ǣ�G��,�����1�Nx�Z��+S��E�ߌT0���9n�7�����#;��`[�6�y@�((T$�l腻��ӿ絳0�(<߇��cHz,BK��T�7:������>��zG�A�+M߉�ZЖ��1�(�c��Eͪ���/kn���@�PO�[=J�2g6��b�Q��c�VD���Z�"qAЭzɦj�K�}h}�+�;��E+(:
�M�Z�pr�X�!anQh�Ј�5'4	��7�?X4�v�!E����qA�)C��g?�ƶݖ?i'������`R��Ê-� ����$�3=�J�U��Mgճ1�j�eV��wA&����S[Zxq�*²����Ά<?7 �����M4It�^@��[$0��$����v��m؍+�)�H���o{2��
��Gκ�"ŗ� NHJ�x�
3�z�L���Ë.;�n����h�U��Im�<L��y�O���Q#+ʀ�H�;V���c��ț�AK� �v�A����h�	�5�����!��A�C((,�f�'�IUh�!�HX(_7'�B�RS�z�؎�a�B��}[{�K_��T��{m|��c(Jk @w �O�	�� U�tUQ�u�!��K�D�+�aDP��/?
��'#BnT��j�E�!IUg|���HD�s��$�Ҥy���ay!y2�O�+�F�C�'��:6���Vj	j��:;���Gg�G�fțY"�6o���ӯ:7U��nHa%���0��z1s���wn�S}*�e��g_�g��劳����rc���?(��졲���N��b�j�`�?�^V��S�d#}�Ŗ;S�?��H����}�|���j*����"-bւ6�<Ƅ��1���w�y�PV1Z	�#���
n���gQ��r%����f��������ɽ�E��O.1r�!ېo���%�����+ό�L3/D��l�
��Yx�j� �P�^�ӑ�(��nv3� ݠ!e��F��8�~�3�O"�Ä�uf�����kDEh�h��9����.�����zί��(U����d-�Љ0HY�._���Zwk�E���⡺>/�w�����Bn��۴\�)A�-��m*EE�w��͓Ӈ���bGp���<�~�Q�V���R�v�d����n��[�蚁�D���MSo��� ����i"<�}�_����S���7��zX�B�*�&޾w���FNd��8�B�Ծ��;���2�R��3^�d�]���^�n�.�c"X��K���ö����s�2ӧ�����\�8,�X�xȪ-��L�+���D�(&%�,��������6���[^��ͬWveL��7��E��n�1I�J*�s۹C|�B���nC��Uv+��c�3�����&�,l:���r�_��q����a�����M`�'�pLj ���B�U9��7ʅr,_I����:�8��������ؒ�A�]R������G��a��[ו7�7Xm����0{�4��z�A�@d�_y�ĉh��6��q�V}�j�� :����<���n���X��w4º�|����V�)�Fey���{��$Ś��H'��Oq��m3�e�ϊ�\:Vt� %�B+�7�T10O@q���3\-�[��������$�1��%��q=uy�D�#��B�
�gb�'_~3�υxI>�3w��d}�<+	
�s�De�E0��g��%?N�ij5C�87Q���(} ��C�WBi��~��ta�>����!A�\v�S�M�y�&�4����8�G�md��q��r�F{�*kw8�H��!߆P����O�� I��^�Ѩ�T�p�8�>�xt3&=3�����L!V3F�o��?�D�ʢ��jQ<��ǤY�U+	��q�+74����y}^�T������\.��Mh��ɶp�R�4_#�8��y�i�2��K�g�S ���@ ����IV��,f�ROm�j� ���CA� �e�F�B�ye��I(@[ۖ0�_�ze���B����x�6��gw׵-i�,���蕋y� �=Y0v[h��Ճ7��.zT��`���>N9��ߝ���w�bO��A�kl%�Y�Ƭ�ǹ�~�-ԯ�Q^^a�}SI�N������g��	����}F��苀��7j�Q>�d��V������s��d߹�K *OQ�6�RUJ�
w$���2x�{o+�ؐ��Z�[���k�5��"{�)�����h^}<�� ��%�1<�|�X��% I.U��c���]�P��.[��h�i�J���t��M!gMm' �_���e�7���ӡ����M��±g��ԩ:+*��6��cwYͽ�C�&
��X��$�/�ͱ�iǋY�D��B����$��/"q���#t]Xhr�h��B��F��?¦��7���%��VW�V�fw�a�Φ�������!k'�����쓐����fzP�E=!:�f�ʻd!q����t|��`"��[��H�/x~��?- ����	����3-����$�)P���Fs�������H�Y�������H-�<�T��{�n\�i}��4@�4v-�̕�=�;e(��B���>�@L�#Hm������3���"�'m��Z�����c� �>}{�]�j�8��(�nm�7E��Xvnoޱ�JHP��6Q��V@sk���͵^��Us݅en����ٔ�s�a��s|$�.��K����ƾ��F���ɯ2WqpR���O�0��>�X��/v ��3��dX�9eAƮ���QQ:oK��R|,al�A��_[.��!���`����t�и!&��%��B�휝V��JL�ͷ��I�Q�/��瞘��DǶ8}N-X�6XϏ"G[�P��9,����R/�7���j��Key�Ge���rZ�G�����_hP|W��
=�[j���������k�4��;5�ޠ���+��0Nz[$��&��i�N�KL�&^?��Pѐ�
p��q}jc��W�<��+}.��x���i8(�o���f?2l�
�'<��E)��$�f���K��:��K�7`���kW����,q�L��VLtl�������� �t�9<ð�y~����,�N�o�p�Eظ�K����Q�~����8�����1��u�LqJ�]=���Q��Ǻ�5��`���'W�����煚(��QN��@UT
��+wkp^rU�<~g�P;�O�u
��,��(�ҲHqpX�r�h��:)���X�>8H���<�����0e�c̦��+ָ�}r ��>��+�澐K�%V�CC�;#E���췭ͳԁ��h9��7煤'i2Hf��e������v٬Nr�ᛀ�sY��N�ϸz@bP����!c�0�H��$���Bm*G��W����d�EO��A��U����e�>���(�C{߻�g��YePF�`��n뺉�ڊ^�h3_���7iF�%� K���z������v
���(�*�
r����겆2	���KRj>�R`҃Vk	Ƃ��,΄sy��9�����\&)v{(|U	A�KKz$��v	��>���)(���)�ϫ�v�ݛ9H����~�"�81�8]X��(r���M�0w �N�Ԝ�P��O�IݦW�^���B��,k�9���+J*	�3H���t��o�lp�D%�tB�v.L�80�l�O��t��T�]�{ڋ��U�i�Lq��O�,���!O_�Օ�!�đV &Q=I�H�A7���	�:��YPa�)���[ ew�����;m��Vqbp/n��h�[��Ή�P&��p���ľ�zJ�v%��Fl���_�&Ŀ��q��+#»M�5�F�{�9�4*T�f����,�<�Y�]�jaa��b~��OZJ�����O���s���ucԖ�̖V?$U�����>�����U`%��I�8�2q��N� �QY��lao�A>P1fT<�ɻY�7��b�w���cz�v�ކ����+��J���e����$d�9걌l��GP$)%LN:Jn��I�f��U�}Q$�$���)^�)������?wҼ��:(�d�"e#�3������ �����8,4�^2�EU��J�6�������"KO|�n�l�1��.�6g�Y���bcf)��g��O��qf�����])���@E�UT�:�G�grˈ�c�Ԯk �+iFQmc� *��l�W>���iXy�fJ@g�m:*��;#��"m/Pri�0[�v�e {]*5�X�/�i�2�e������OG5��,+�o��F�j�F�\����W�Χ�.4����3�(�M��-�롾<�����M���!�{�`xGr*Vɾ-�G80�{���ȿH%|x���>��:�|�撒�Bz L��E�x>]�N;��Ԕ�������F��tt\:�.�8��B�Hw�*Ϗ)z��u.���x!xr���+ ��6�3�ϝh+U!�YlM��i�j�������vn�I�R������)��?7T���>��-�]��GZ�s}<@O�����̿�o-����nL
B��hw
�1$z�U:�����L�-hȅd�:z5��'U(�O|<�B.��6H[�T��i2��V���`�[���*�-GLS+~&����q(�[�>~!n�^���4��a&�|t:|O$y!q-�n�	�Ŧ���0 n�)�MN�W�lKD}�	��G��
��wr�B���p^��ȆH��?"��'6|��|��C���B�}u�e=]�jiR B
yP3�.�É��㠁LI@�kvv!�a��:h�ԇY&b2�H觠"�ԑ��^� �(�(���.�)7�b"A��n���h��0L��)rYc�̱
>�|�'*��ax�s�Tp�sF�9��Y�'�rc�o��̲𯼙~��ӷ\oG>���z����6-���e۝�h*T}�Jx�l�ʶ7�Z*��k��ANsWxU��Ln�tB�M��S|6S�h��W��� [0�G�B/�ȨW[y�\7k�I,)�蟐���.w쓏��M���e R�;)X��9d�J�X�4!#Et�&�(�*&}ѫ��)�ng~�SE����m�Do>b��l[�y�!ؾ�0��(��<q�B�ݼP�Y�����ꞖD5��FHDM�rA`JD��{&�:8!W3a����P����j�o')��{<E��f}P����N�xq��c�,�V1R~�0�IrR�57�Ή5i׹B�LH�D�e�^�ñ�C�t�c�����(�*>������J+#��D>8�!�\�=b�}�G"�jun���6+X��!���%��w�l�u��{ �������6p&h��ms$��;��C<1�;ˆK ��c���S�o6��(�#�r�0ٌ'�si�R7'�w��<���:&��)	;�-j���x �y~�:�����:�V[M����/Xj��z��-��B"�ܨ��E�۲?j�&��,�];����Х��#YQ)T�A�z�[`k��/ߜLx��/G������4��#�}AN!��GQ:-�9�	�֝�bw�>���a~���z]����i