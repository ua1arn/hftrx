��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�E�Է��� s4v;�7]XЖPMٺ��6:� KdR�t>}ԑ��z=�kx�֫�
|"��V�~ʎ�xP����7$V8X3B��'8�Z��Gv���[�`Lg�L�Kno��r��������Q8�	my�ۏq�.�n�������n��&���x�W�kˌ����&p�^��sj�ۘ$�}A� �S�vә�vR��� �0o��F��zb���"0�Ph�5��:`^�9��qy����F4�X���S���+f�> ��Hx�n�%=�C;�m�igO
셝-!�a�'%,�~p��Z((��O�5-ve���)V��/ބQ`.�m��<.�ղo�Z��5V{�@S�����{�����1�����DZo�w=���q�PJd�x�ۀMB2������@�mkT�u�F� �l�6��'�
��ԧ���i+��ۑR�)�f��h��֬�����HQ�*m���y��D���ܣ�#U�t��^��u�7PTNXZ�[�#
�T�)K�^!��~S������~N/��]��p>��l��c} ���?U��E7��m�W�I���R������m�#d�=n 
C["��ӟ��_��;�nWN~��
�-[>r޲O7����7������f!���V�j2S@l*>�g�GZl`{�EMx�	���". �T��١1�"��[B�p�i����Q  �v���=|p5W����+O���Jc����I:�|�
Ny���4�7�c 9�*U<<���+M�6O@ԓ+긁Ww6��x�!:�����ʌ+"���&��!\^9>?�(�g��=YK��7LmjBft
bF(�o݄$ʑ`���Z[ꤽ�l�F�q6:eH:e����ε+jiDȉL{�ڡ�^]EB�C��w�|��>���\P_2�ǡ���B"��w���i��+Ɨ��kd'����)���
�'i�C�S���K��,���0܁��m��y֚�B���Z�	Aa�=Z'�F[� p$�bi"/"G���o�Fr��z�a�/�i�X���f�P�-%t�n�\��L1M5*?�Y�gm�ҹ *-�ۙ�$����
VO�?@K|�o`{aG� ڎ�}X݉�Vh�l<��G�����A�Ŷ�DHT8�|�>���TOjƓ�Vm�i�C1	}�!C1i,�<A E�(��:*�!zj��K{�g�י(R)z->=l�l㣥�@�G���� �]Ʒ��<w�%8먃9���j�)�9�6�` $��jr��DX��ԣ2l\��&�Vm��A��O�<#JN<��R����Z�x�[P��0��%���#!8�����xqK��!��$(v:Ĺߪ�%�8=�>�Ew'���'�����
�2~��@�~Ou�����#��ZPN��Z�@�����\K�&9[����*�o���]��h�2�u�����ߠ�^-������̛�ng����= <̂�ş�$���(��c��@��9��I��6?�-M�&ECV�OKaw�I�x�Q~�.��0���'N觊���_4�:��-��--�t0��]���Q_����NK��W2�/¸ֿ8=����|��t�4�aWwh��vx�K	8Juo!�f\�ȷؒ�����̘Sv?��AP�Td��2�-��ƣ��EHl��:�c�@̭{�ϰDe��1��cP� ���\�i���]۹@}9�᎔-6 ����1K1$�� ��g�'<��.O�M��� ����0��Bj'�.#��
�A���=�s*�;���w�Yk��f֑f�2w�e˞��C���:#�i��]-���R�S��U��}QA$�T!/�뙇d�P��d��Sj��O�u|f�{�C>F��ĩ4$M"EU��{<�UN�hC�0��X��$l�� `�2�-7�z�>vc�&�(�ir��s�|�-~�����1W�1W��'��z��A��`k ʳ��'�U����>�-d�0F\�W?+=\}L� P9�"jk�?2De��ډ(��k�������Yr�L ���5Б&m'��6��I�,[\�S��p���m��8��S�D�S�t��#R�sL�W�[�F0�%�v�SbV��%f�X���s:Yj��@������h�lXH�	i��>��֘�әh�-���?�]���y�+1���4�Zuz�r?�ڪ2�p��D%����ƿ�8�轹�I%1sC��W��d`o��!�pَw}񍩞Eod��E�/I��6��0w��La���c���R��WĒ ���+]l��Qz�tD�.ڤ�"WҜC�sH��(�J�8��v�	q�i���%�ՒI���|>�(�Ә�f  z>d�h�]'|@J�+����upjy�%!a%�A�;��*<4������� �G�vt���5]nxeb��:�&�%2K2a�x�"��v)q��J��s���M�G�>9�����g����T`�vNy��v����4�!f^!=~�5�E(�����6�^v)��rΦ�t�lO����4K[8�p�U�`o+�I�	�ZR�9��g�(�l�B|��ց_��_jA�r���r̬�f�(ee�����S�~���_T�ª�d�����������}�N��3�C��WB(_���uݾ����`T�2�(��\�"f_T	��D�H��	����dۄ"��R��yd�����ɏ���3�0�c+&5��g��S#���K����6B35��úD����0�.o�1_���$��\�0�ߍBQ/�3İ����}�K����|U#Y�8�Jt���H�� s�4�?F��>��Z��� i���2,@�t�*҃Y��>����uS}��SI|Z� Hzȼ��#z������*����˥_���>�o�@�h��4jWt�iU)q���k�\�ˈ��y!@�H uɦkM�8��s�閡���~S ��&}�5(3�Z2�a��4�m���2@��&<�tM,0**�_=�����qB�G������~CƖ�=���&�&V��|�Ҧ����y��>�DP�rB��8f�b������G�ale��E:^����f[��:�=�č��I���ds��[y�"W��0E5,� ��'��M+�n�h�9�c��&� ���X~v���]�u`:@��b�&%���ǰz>c���4�������1p���6s&��AWe�L��$��f��$z�a��