��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7�ь&t����l�e������as��U��p���t��|��=�<�4ХC��-<?_a���}B<�͡��zaRX�oD��I�=�Jz�'���rt
o�G���ֿ}�\���˘�`���P��D/F'���mZ�:������Bhs{
��-���������|rJN���ֳ��]�����-q��Ip���¯���e���'C�Y]�ٹ��@��B@@���	2��,�b��.���^�n~�v�N� �=�b,�ƅ��c�qhCw�����Gwuc��?�ۢ�6��.ㅅ�Q��vq�M����}���ٛV�U_�gi�����-��'i9Y��g��So���>U���}ۦ"e%d��u��,�*�kD,�+|�_K��{��b>��b�˧�Q�d{Ss��o�@�3Ն�;ŠR���E��Nb�'��eĞ��ge�G!�p��Xأ BR���(�e���tA�-�C�`���.E:R�k�NdqFs�ZC��@�0��U����3"��*�d�,�%҂��#�#{⤆l��?Y#6����~��}�jY��N�����B�l��l�� `s��Ëu�B���������Z�L�6�DyymK������l��q��ؘ���M�I�ꂱ�8=���ǀ�]��oy����{d�E ��F��)����R�$GNպP��\(�'�_M$��yy��*�ε��e���གྷ2
s��.���G��#r�͏���4���Q�îp���V�R��Ņ���P���v���U�����š������q�Lw�DM�.�}��n����>`�`	��7C����	5w_�A�'0J}��)�X[v��,Y�������)M�z��86�P&�F� �B����wC2mʄ�!c;�k�����"�'p��9N�ف�K7�v����*�e9�)'��"����ɯ&7"�#�15겼����=�/��O���݁l?��M�%��=��$|��y�(��ٿHW���\l<���,���]�� ��^��<߃p(N\?@�g���Cqp&֑���@'������W�Leb�A�OFfҗ��C41Sތ�>���nk���G��L��ø<���U�l���i�:e%cl<ִ��yy�t��E~5vͶ��u�d�R'���V�d�H,S#��%�$�Ȕ/T׵T�]�y�2kqt�{�1�o3/�/��s�ս��7�6�VM��l#^}�oy��|����f�)_���,��$n1]�FU	h+������P;`P{�"�*Rg�m������D�P�X�g�[��)f�RwLSـi�~�F��4{�	r/cfx��5!O(�����OMj����{wUU_B2}��Q��[���!S����ϴ�����Ê��ќ�+���MJ?{2t�L�s�5p��:)����!�_v8;c�cx����c�7v�>+w�7lY�EaZ����c�͠Ւ��R��Y�r?ӈ�[� �T�j-��?���#v��"%w5��Y.;�tă���V��c"̭-q&����2U�o�<�"k9���0r����y�:x8�e�c��9������������s�`��op
��~g}��n2kUBTw�H�H�m�����jc>3�=2���A�V��@1�Hmd���� P�"D-#-���ʥn�$��.�W����J����]{�!$N	�+B�g������ĸ�������a�''�ku��_)'�S"ÐP.�<_A���r��%�q���ë!IL����rN� W��f �1�������a	��u�0>�1Av�B"��_�u�P��X���� ��x��cs3�I��w(h���om�fCf0�Q#6��Y2�CD>]4.���H�>�!Lz��ػBJ���!3*��:���U��~1#�ܧ��C���aIKGR	�b��5
n��9�u.�к&*�.�.�m�)���Ňm$���c�fo����yM0�&���s������!��Ӄ�8�����ʵ�q���erKL&mr�R�q�\¬k��s��RV,��g��zo	��ݐaG���k���p�q�9x������E�	ٓݷ�o \���jxB�G"�T���=Bm�w���P�U�x�!��QGw���7',�r���r�bM���%�k �.�Hއ���	�xc#�(�Vk����(���E
K�$��Qw}�1c���<�H0DP�T�V�AV��+��' �y�[�;���L���:��i�ntG�I�cNd�N��Hx��^ChXM��)cQK�����Li��$z@n�}P\���� u�0B �Qn�)��`8*�J���S�ٝ�^�`�q�I쫶���%;^i�Ϻ���u�4]<����|�
��d,��K��(-h{���y�C���H���^�3u��l�3R���'�Y���*bj�)����y q���
�\b��Q�x��C8&�z�{�(�^b�:�g�h���_����i�7T�d�_�XEFo4\���Ώ�kq'�A������{��w@Ʃ����<**�;%�Q!:�D���=&����/B�(���^�����Qi���1l� ����tZ�bs��:,�a���<��P/�w	F�@�,Ϧ}gI�x�0B����b^K�x�$���n١?�N����;u�x��F�Ad��d��h9r���e��hL=<�޽7�������Q���pm�t��H��	�O)���+������g*��V%i�-���,��<]	}o#\"�ZO�^��'}�ӝ�Q�0�c�/gxWǎ/�Q�1������@����@�q<��������W,�jet��/`Q�i����2�d��3�d�`�����M�-�e�3&���o�mS�K��iIOV�|N�_���N��8ܵ�J��K��q-��.������-�%���p����J�d4�?�\ʬ�&p.ճ0�a^���&�^@n��q���aVG�Ե#*�DG){��'ً���N��T�^]��.�峙���ᲆ&�$����v��>�1	�#Vl��:u[�����%���H���Q�p^w��l���P�� �)���$�s���H9w��4s�_��YM<P����g�F�F�:路y��$7���LetNk��%ڴ�m%_���n��6�	��\�i�>F�V� �=Lc��y^n��v8�� �Y�|���Q[�b��50l ����q"{`-Ma����)
v%"�=;/�e#������J¨h�@������#c�xX����O���V�o8���*����4�L:n!~WWd�_�r�EL�+YH�_�&&�����{M:QCk�=T�B݈C�8w�w	hD�|>�)�� c�}W��ຜc��i$�M��K~�оY+=�9O,k!:��o��V���$���Ȇ��x����ϑV4�����
q��"�*^���؂t�j������wxDY康Σsț��ڣFH_�	s��|��%��H^�tu��GqX����G��L�G@sE���Me�r�}�o�If������ Z��/d8�*�ؒl���7=
�,Z�,�Bc��Md���;zK
�ꎈ�e/�Jl�SR�&����[������^����M�lR^���0 �?�%."���|�n�8���Eg��p����h#���^��-X��A�L%I�܅M(C���H�=<f#q��#|"���ǧ�pt�Ӯ��Ǯ4��(��䰞���
&E�d����\v������z����m?M�n�ғaf@O���3P��a��ّ}�רb��_CU��Ke:b�XL(K��w<������W�����|��s[���h{yy6]R���t�=�!9����"��7�-�c��N�������R+O��9vYX�.2��"1Zk�Yk3qZ5����g�0�߮��������U�k��~�	�v��̿�k��U��)��]��7?����	bM��g�a��SC��<$��	����}�R�@G���(ge���)u]����X��&���֧?CŘ�������)�z�W?�W`�Ȗ�m������u=K�A6r�p5�D�+�;��+-��'�K+#w��.M���^b����7�5���T�i��`�h�2	r_�+��65���>J���P� ��o8=��W7�m d�AT�Ɗ-�����^#ɣ�����0��\���
�}X�����U��2�K=Nb�!����E��APgz&p���@�Jr�r�e
F�,��"r�S
p͓zlT��۬��ri�z�U�R�)Rk1Q�j���>���a:�ilĂ��St�+q�%ˠ��q�X����u��7�^�_<vPW�?��&��YA@���:|��|����_�Eun^��ꌦ�p������YYr�㺾�J%��XgF�� ���������s�-�F�l��6�h�ކPˮh@�K��S�����0'������i�NaOW&=�}z��v��q�C��#]T'H�Ix�5�t辐�>8p�Ϯ|��'�4�dF)��٭����Ka��Ei�X9��@W`fb�B�Z�+�g�
8��)J���b����D�S�z.���J�)���4f1H<%[���O�]���x'h��T��f��'��7YD�, ��Ƽ[�F����N"�FG���bY���e�^���@�c�1�=��懶��%J��̪L�����k�Q���f���NY�H6�F���~��3���X/�>��#h
��Y�#e�N( ^ X9���51�	\z|&�מ�pM�2�N���<+�s��bk�c�r����i�#�B�>�km���t�Nrj:�7ZoG3���8'#������ !�=��@���E�I|�E�u�@�125"Ir'*���^��x�S2�mJ,�X%�"љU|�/�s�����w���h�Ҙ�L7�x��E b/��4�+���4�G�P�Ю׺�WF��w�L0Hf`��c��uۼ�i�4Vq�%��jv��Z8�QO?@�@o��N<烷&"�:��T�D�w�s��tܲ��i3	xKP��i�(cHbGTfq~!�=._I�X[ }I�J+>�;�'�#p_�O'CL��x��B��򅘘���x=�xN	�}��D���ʀ���8���!��q����G,�A�'M����y�%����F+�a}��$|��Qq ��OZ�bEp��1���R8{�Q��R?���܎��c�2{%oYdҿ�T�l�W�{���E�
�q�ڝ��3���lk�Æc',z�xy�?ŗ���UR~˴Q\d�AA��7Jv����=_��K6����@E6������s|�D��G=S��l�v�r<�$Si�����7�d��y�K>L��������} .$S%D����pιL�����&4���?h�l�Y��jA�4�g��[�ݬ�StnD�_NCm8�(d��@柄tó����s����L�AL`���L6���NA��	!
\ک��.�����_��z��>���195�̹YU��Rs2��Y�ۦ[��p�������X�{���D���j��>1	eb�D5���x?�7�5��N ��wi�&�;	S!$�I�k�����^�Q���bJ�I�)�*u�2\��_qz���N�.�|8��#7m�	1�������!ۻn�zMp(��3;�թ�`�{���A7��W�ΟZ��V9�5'��D���)<E�@%(����kn��yQ���� �SNw���4�,���d�bOgښ�M���,2���$I����g�ڕ�$�K��OX��~��`�a˅%@��� _�IDB�h��������A�b�1���~�Z�	^�d?	���TyqB#�=��?���	�G@��g�(\����`_/��hM��o�߹�?�%W���<�_f��Ikc>�wE�g������]��G���F�����F�uC��8hX�N��>��T�� ���&�6�a�w��=��p����r ���Ƿq�4���q�?NPl2�gÕT�8��SIF!=��Q��.�j�U���|�:7�Jt�Wt1>Et����?7��i"��]�d�>vshš�=��������@������Z�WЮ>vk�§*}��<��������,ae�T�/�Ϋ���>v�;U�PӖd�r��Q�k6�� �M�>5wZ.ۖ�0g�[Dx)Iہ"�'{�.Q�	�=Qz�-x	S�k�п���8Fֶh+����A\���S����"��44�Ud��WEbj/��k�J��������QG���xp3]�?�K�_�|L�K�H`���Wx��E\����>��ѭ#PY�L��R�:�;^�Y�ؔ�]�W�qy�~�e��|��h�`��|�/-'J�_�X�����Un,(��B�Qj,Z�z
Y��1޵E�
��E���gCoF�e�hY�mHt��	c%uz�=Y��%QZ�yx�*�c��j���
O~{�]2�^�)۶2F��%���C�E��������M�S˛���qa�fj6�a#x༿�k����� ��V���+��=d���� ��X.n���f4��X�@��'�R�����6�iM_� ��~+�feʄ��+��:������SY�P_��{ѨX0�lFL�E\̞1��Ly��-y(h����lL*��^��MmE�X‪�N��'��d���H��ˮ�`�3��,����9�Fā8����2�Q��v�m�����!�w���aC{Ʀ��:�GBl{��D��+��\���tQ`�p~n���Z]���Z��p�[D׬������HWNAX���yK���6&�Z�ZٓnC���$-�+�|Bš�di���!�<l��ׅ�S���������5j�-A���8�I�F�+���!�.�
ڒ�Y9�xU�1fhTxh�	ɺb-�$P��k�	�P��j�"���l��=��.��}.|R��>�����ǝR�+�k�-E���V�0U�TO�
$8z�ܳ�������||}yǔz�){��u|YCN�d7�*�}�1nk��>Q�Ã�m=�r|Vz�%�#�8�Ix��A�=�f�s0�
�\=��d��Kb�+���5� Yl42�o:{��
w����2��No�m*��w�9���*p�g2�t�7
��X�e�z����H�X������`"<��¨�2�q��5���N�ͮF����q
�