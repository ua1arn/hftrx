��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga���<�\��J�ιϛ��u�̶e��I(�LJ`k�)��F�Ϗ^�a	X�86�|�tb^,4TVb�y�I��}(��ΙQH��y}
�b��r�A9�S�ڈ�&;${m����o�F��`��oo�"���{Q��L�>�=� ��y�������Z=������� �'�����晁�Wu�T�)[��%g��"N囵����:�}?�Ña�bm�����)�6/o���#�I���8�aD��g;��E�sۼ �ĸw&�M�hx���~�Y�4�,��6�޹��~F�Ӟg<p����g;���Os��*%��)�.<++��XR>��#lY�z��3���<am,�ٚ ������|���݁�K�����Kd������˔��S�ldw���ʜr֨���`��%p'�.N�J/2�_&4�J���3S��#���us�N�I�e�~����4.}���%���5Rh��\x������5>�$|�֘�Y�$ɬY�A0�2�9`|����R!�L���1䫇��q���h_Xӓ��S2t�M�7�f~ !�>9s�4�{�/*E�?�W{A%�ph���0Ԃ����b7T5���#�=��������!$5�H6J�O�t�&����h���7���s�w���iI�}||ْm��}��"����s�M����ٵG�����>��ȉ�*����MH��l6+}n��]q����^��K�V�o�n��w�/	?FĴ�9�**	���Z���i$ ��Sm/��L�\��p�\�X5W���'ZVL�)<��	����[��k��u���ҙ>$���|�.�u�Kuk���^��k7���ᲆ�����S���D���϶MUf��_����~Lx���(�����#�TWl�F��T������W��m���`����N��_�r(!�_j�~�2���S���?O���&�gȖ����i%�B%��/W�������U�> WV���^���X
�#�M`Y&���E��[jlWDdek��Rq�T�f���͵V�K���&nAc����I�)��v�č���������JXB�Vv�zs��Nr
B�o3p?ڋ��L�3�~�-͟H�ug�~;On�n��#���Y@͙�E���Jd��h�g��Qw���-����gw_�;���n1G3���t� ���#��D���K�9޾>����\vA� ̬I����@�"��Z��P���z_ܸܴ4�3{�,T��-��Fp�EC��yj1~�����t�B���gZ��� �"tb��}8�&��HQ��P�.���4 �b����2�4��4�j_��loD� `)�L�-�͠��/��+N�.��y�n���ʮ|�$�0r`�^�=�̼�_��{FZ0�7��E~���¼��8�����_*lxM��5%��j��h�($��ׅ`�ˑ��:�%�={�k�N�XY؟gW0�z)�F^m�e�Þ��a�=����D�m-{WXB��HE�+?b����L�I�ڳf���eVb���x�� ��tV�N��JKM��d�����o?�=�Xk��+Fo(�'U�~�xu�͓18��H��-�ȟ�|P��n�_G=�慤���_R:�	7^R�d���[ i��ʠc�0��x(��3e���l����S�� �U��e���`7����5vv�`���G\x_#�Am���H&�e��k$x��U�el���%�o],,p_�@[��5�<�9j!�}B��#�{Ѥ~_�VoBd�Zޑ�[U-�E��Q�(�;��g��~$��=�v�w �SC�R~�쨶��1*�{l1x��<�	 �b@;J�N7aS{��Hr����a���G0p��]l_! �뮌���%���=�U:���t�O�e��r�I���Cd�ǯ=7��I���p�!�i03��xM���u�Jy��2>��8Lm8��k�&��S���Ϻ`i���q� �J`�SU�E�b����g��S��ԡ7U���t��@8pU~����:T��1�*r�$���x^�#e���C�	Pr���;���Xr�T8Fd�p�ҷ� D�J���ۅ�bº�%��B�U��ک��x�Re�圆=�[��o��I+H�ŷ�}�Z�m�+��h�[/3�uxӘ�[W�_��K��)Z=�Q�����z��w0;ca X��vG�͝�ȣ�D�jm���2B �;'���R*�f���'h[.bw��e�Q�=MW�h��=��&�
e�
�FX���(R��1����_���D�+��TX-�$Z1��p?�r~2'�˶0�rq�mS�9��%v�_u��~��+��A���+0�!+�9}�T���f!\��ِ"�wN�$�n��$y�Kz�,.�'�A�U��<(��I�`����C�J���r��q+��;�$1A�#�M#�����ur��RC��dG�*��"C�0uo����D[.����)������~"��}u�ޠ��x��k5�kSHf"ɀ�m�Ͱk�5�ܴ�J��������3��@����jao�)��JD��)V���� ��X"���5U��c����}��;=�&��sRZ��9ͺ捃���b�L]>�N8%����4�a9ɾ�(�{�I��4̓p�z�eXЏbEj]#�\�k�Fڷ]!MĦ����8�쌂��v�WQ�(�~�]�d�~g� Z)4��4	�����*��U�D]����������+C ދFp���Q�������^i�ǡ`���2�$��(T��]n3��f�MAQ/��A(y?�$wU�S:Nb�����L���������*H�n#Sӟo}�z����ʌ�'�Y�*�֎��b�}�����6wq0��,%�[M[&�6�;�Cm�N���">S�"�Y�e��U�m�^;�`6/K�6�pU�Dh�7�i�#1Ar{udY�Դ%����F��~=���$>��pq��e��kq m��~[F�iձ��Lw~ݤ��Q�5��-55��?pE#N@��(�ɇ�^Pi���]���Z�/o�������:zr�����Q�Ż����a4y$7����͙�$���%����)¬��oI<ҹ��1/��C����#�ǏZ�v�������	��^�:kI��g���a�<�ŗ��dj�(��'���X��<KwaJ�dV�ϸ�ܿ����(�b�0��s�.a>�k;qWq:(Xn���LM�A2O{�0�	X`%g[�������l�ҽ&]s	��Ő̑�h�`EU���V�����J��)T��O �1������p��֓[yz5l��&:>�P�'��J�0V��,e�b)A�!0�QM��Uڳ�4�ump�ye�Sd�����Z����u��ak7* ����O����k��C{�u�΂"L��|)���,
�3�JS��Tz_�@��.!�c�w#O��Go(X�R�#u:"�+� �q.�}Y���M�T�J�Ӕ�ISl;���t�d�Ʉ�#��[�;Ƀ�Fv7�
� �&��p�3�=���С"j�������[٫���[��<p�ʷ��z�z$j�xR�hR�8!�P��X�`z�@���^�\��b5�:Z>��A���bx}�!��c7���De�M���d�ۢ�\o��Lp���>J+��3�˒�$��''�i�#A-���I�_?�/�&���@�G��h!��bs���e!(qM������A.��@��L�&�D�+�	��Ȥ��4p_�~����S�/����e}��7��N�Q���J��mI�_My�n�u��"F���1|�� Kě��d������[�[�AӮ��\_cyܛa���Pt���r�`��!%�҈f��ZSо}�iy^pT�����	�!�WUmPEt�lZ�͛�g�e}��pTN�6[i(�w�qx�}�A���Kԏ����� �px1�l���ֵPc!91�9S���%���ʵ�?���g����:�Uy�V�՚Sڕ�����t�V:��R�wZc�M1����� � ���Ͷ��lx��붴��	�������}���v����.��Cd��>W��3:s�&�_�JO.�GTG����N�+�r�T� ��V@�X���Hʇ8��e�hH}����+�#ScB���z�E����he6���, H��Ǘ �L�8��yEi�=��	Z�����b�@��"�x�!g���Es� ��v��@��7�AT3�"�2o�pt��U����q��b�i q��.׈P�2?	�h��fO�L[0�U�ZG�kjMYN`N�E���;���ؖ��K
' ���q�����xC~u,�U�>P4j��� R�v��L��v�ɫ�PC��-�߭����57'�ʘ\��}��>���S\x��8�0��%I���/3&��@��'/��a��3�r�˳?}z�H�ؿe�2��� ?&i���uм0�����:-��2�^|���F'��]�^OI=Cl������ ]�^]�Ǭ=�Y��z1�CU���^�KHgd<�WX26���䵒�B���������A"�WM�hԭM����T^V8]��ޗ�����i�9����,0ڌ��������f�����$�rm�7�d�Й⒅ވ"ţ�2�L���m$�h�c�����[�)�Б{֬���q��� I����}�1�h�B�BbS�Ƕ\L�i�Zi����0�Ŋq����2uS)_c)u�{�G�� �@�
�a�����>H��O��0H��f7C?h�{��$��UyW�5��!�F�I���O����T���lt6]1�y�`� 5�`؅�6��Fe�>ƅA3�Z�d?��+��ʹ��U� !kPt�|�~�^��Bb�b(��{��1-"�*_��cf=��<[���ˮ1�����Ef�>���(�ӷs�^�,�A��Zr�w #�G��+�o`j�qH��
� ��#�.�"=��� JE�0�(���m�����s�f&�z��3�ܨ��V���Q-å% ���	~�0E`<W�^)�<�qG,�K㎛3�E`=��/����*8q�]?XM�ů�
���υ��b6���kBa*;�?#/lYԥ���ߚP��Q���7�CSj�E
��5I��8�th �&��B��m0�pT|X޿D�~
"�Z=�������s��\8�!y�/����gS2�����0C���O�Y�P��斆e�y.�,�?I]c��]��<4�@?���%�_Դj�J�X"(
q	���M|��2_���p�
�1��Ƃ}�%�3e�-+���A�V|�%���Џ�,]L��ƢzGZ����zW�XK��H>��Qכ��R\x�Q|Y�h/S�m��8�@1�q���߉��%��bi�$a��*x����Q�DZ.��fֆyg�E�-��b�>b�����B#�5��w�/�x���p��A����k���<�����!�d�r�zF�6�6�>d~�b�T�ȗB+%��7��_W5���v��ȃ�Հ��n�oL�q�~��� ���0 9FctB��~��A����1L,c?VDyX���=�5,��ެE�6�m.X�<�'2#]�L=��v�NFOL��]�����S7���S
��s]���	J',���"V4ʡ�-s��Q�wWk�0q�y�n87>k�i���'�½�"��> _�ګ�Nn����@�[#�v���u&���/�Q�J���c��f�3I?���!���
E�9���zI�Yja~��tBo���������������ª���))~�[W�!��˘���Q���n{��]�W�����O/V��0ܐmch�-3���q�������Tü+~�4����ZZG��|T���Eny���'J��������{������Ζa�n�v�H��L��$�f����
�8B������np��J��}.�J\�a.��1�5,����fm�TIm�'=w��ʅ�?VW�9�8K̤~h�N OWX�]��)r���#�ݖ�/Gd���nPE�a��<�)zf�[�H+vg�s�,6�'�p7��T��
M��V3-.��J+6.���O>�#F�v��Á�>j_z��;���Lи6a�N6ou�gʶƬ���s�؊E�Q�J���4d̀��no
({��J󘐘M�j�c����ԟ��UM�&�[��������ٌځe�z�B������&�*X0����|c�#���i��V��5\�ѿ�%�^=1�t��3hi�Z�`})w.�@�E��7�����`��o�
��T��;:����=�lmw�4p#P��� J�����e�vڹ�������EW/��	Esb߄�'KH���J��52���@���4-�����R���&�pH�{�>}̀����������K\
�J��a�|4��:A��6<���l�,ІA���_۟�������	X� Qdsd@ [�ͧ�A�'�+ޏz?`�v��Xp�*��Oլ��L)����aF�$��.+I[�]=#la��{��rEm�G��"�/�3&��r=�X
 3k(9����F�����υ�������H�1C� }��ȷ�f/sh_�f�2�x&�w��7m�× ��H1ۥ�����ĥ,�R`�t]�z�Vןq�43��ơ|
_�ۮ��E�rJ�>{�_�~�>K���fY�?2s���p�'�*�,�Y= �H�j��,yd.���	=#w�.�]�����c�-o�'���y��3f�ux( ��4�Gh��|�ͣ�U�Fi��!�er�@2�)t/�!y(�h��ȮC��a�dZ���&�z����=�P؀ZiN*���5uh��ʠ��dڰ/x�[/@��ߌkT����E0����7�e��N�6�/|������v��b����+ H� >����:b����Ax�m�!s����]#���}x_��+N��r� J�J�\�/d8*|��`Q�}=T5l�RXox7�E�q�v":���):k�	`�g�w��!����$�*(�8����򇻇Pf9.����خj��ߐ��?2��]�Ar:�}c�� T�oJX'��JN�ѯZy<���K�l̛��2S4�А|�N��	��Qz�%'����������!�d��&�-f���`g�~�N�{&콑 ����?o��Z�de	O9̋%i��0�縃ŋ���H��t��cY�I�������ʕ�뙝��Z���Jyf��#���8���!MJQ7?Mpu���v	��fHf��km]��H����m�L�(��\��-�����oIKA�R���9h�ŋm��u��o`�mQCh�|�*P ���m���P{PAR6�Fe�fߞ����W��S݉�"<�N��N��ɃZ�����0i3��.ފ�1�����l�U*/���5㹭qG�99�t:k�fqN_�:xD5�������0[�Bby�FQ�d.w�أ?y��'?@>n�?�m���_8�q�������$� ����ѱ��p\B��KӹN����7��ϻ�܅&��޹�O/#�����V�gT�����>�"������n���7>5CE֫�d+gq7FZ=8��]M�!n�h�Z���>̽�B�ETߵ��F)�|��weG[�QÆ��&?��-&�T�S:��R'�")��3�e ���0�[KHaik�E a�en�Fr�Ͼ��R/���A)܇G������ɼ�̬�m�����#�1���[tt 4��ҁF�'-�m~0��h/�t�[�˒�PɌ)5��#�9+V��x�44b�: � 0��p(���Oe	@�a���b8���E�:Tw���Oˢ��y΅k�zT,�c��q�Mu^M�
���[�Q�U�ũC��9��7|D{��O{3 B�ɃӂЗ�i�E��|1c��@;�Mt��
s�cR�u�x&8�yd(v����v�>@g�kT�c�)S�Ƀ�](�s�n�j��/�J��Z�eZ�+C���_�W�]?YONtV��:�bG�ָ��tW��m���:4�������Jl����KKqFV���և���.�m�!����z��Pװ��)�X�tj\��NX-R��f�ֿz�+Iٰ�@ړ6Q�Ft{b��������Y������UM\�����b�,�UQ0V�����SS�p�oP��<��<���Èw{E$�����8��@㗜��J�/����t�r���-Ǉ�f�#8�=G�m�hPw+4	��k�ws|�w-�D��$[}%C�Y�c�6�akQ��uxt0�A%>�So����M�C��ݰ�K�wڢ���NN�c���I�B�l��u���ʎ��H����hI)��
�	-́����#�kPʗ`D������T�Jޙ���t����%9(n\	y��҅������&�8��bng��Xw���	�"�^�:���IG�m���i��g��!q_)Wq�^�h��ɦѦ�ڴ�cr��go=�?6�Պ�(�+��lSu��?��+�����E+����$e�j��T�d(J���بd�Jف�����8Y���o�M�m�U�-����u��Io҈���wj��<��r]�p
�И�Y�错���TǔW]����C�Pեxx���-���d�`�S �����r��.hϜ����M��1�i_+1���Wƅ�0����6wgۚ#7Y
t��a�m�96�x���L�C�1t:�����ΈĮs{��<��氲�*��b��g8���ny���V>���́����>O�^˨_��Z�jU��/�g���Tt���u{��˺��M������2�:��+b��0%��I�g�hEs�'�%f�(�`Ap�B 2ץ���2�#��q`�	��{���}�jm{Ǒd)�h����B`��+���0�V �Ж��p6',��� 	� Q�����������02���B����u�'+��&���]5�B�"VHɗ|g����7@er�~`���'Q;kõK��|C�vip������Y��%�κ��P�;����g)3�;_��a�csޅ�O��*�̀����h
Jn��z���!�6�L�ª�>��X"C	,����z�ȀLdD6������U��3{�bc~~���c���k.C�.K�xS:ŀk�1���� t����R�$r=�1-������@7�{!�C�ے�b�N���M���9J$��4�Z^�مy퀸��.�d�����W��~mۮPt��
kc�O@��[��L�����`���ฦV�3����{"v�ᷩ�	�ฌn��W�c�*�cf��<���&
�Q��
U���cy��W�<�p�U�@PЇ�	�{*�B�$��D��R8��s|�q�k,��)_b~O)���c'�|��p!�����"��ۭ�8?��BNE;��1X����-�*?�SU~�;��F�����K����
P.3�h28�)���3�����Sx���E=;����
�X*�`��ݎ��=���l뒮i��(p#pɭP(�Q+��(-]yz	�6
j�=��������.G�z���6@�d�D�#�g�q���ǘ>`�*9��l��
���Iܳ�V�W<۠���^��L�G5X~���;FP�"�8���?��v�[���+fC-r���9�|��I��u�[��Nu"�p�ء4|�$=�S��G���A�
��ؕq&�����f�Rh�����߳�{F`��u�����^[9n+�8�����P�������2�#��S�ܜj4ʋ��6�_���6�b�t.�&�'M����A?�����H$~�Ǎ&zs�ߑ�.I�9mKg�0�4И� �:���BpרH�,�\�� �.h�Kq�M��`r��~H��P�<\�ȷ@Mo�P~܀�DR_v}�j��b��T���7=ؽ0����˦s�������>�1I�?����!�f�A��U�@f��z?��j��J�����0Z�c�~����A\VB⡄�ߨ�̞_5���_LH~V�LzHta���e����;
��<M�|����<��X�QP6^V/��k�5+'@�� ���� �C�p�H(ܢy-!M54Sjq�a����T�ʰ�l��w:c��v�=����
�3;��B�G~��@�ݼ�kE��_{�k�'f\6���.N�G�,�{�<�ڄ3��e�	e_fd����̡�P[|��˫gm-�r��l�0x2���`:,���ۧ�S����ef�&5��ܞ�Y�|�FS���Z'PK0�{%��6F��A��7iFr{������1g��}?�haB�Z-���bP�L#UR�p�Yƻ��O�����-Q&�����b�}4"�A���ڕ�9���C���1Js�O1(P��V
s�x���e�r��r�k�Wv�&W��$s֬��c�� ��ђht��v3�JQ���дp1D�)ի����J<݋���ˑm���%t爟���U$0��˨�H���Q�ҥx!�x����ۀqS�nx�HP���_��T�[��W;�W 8�B9оҹ&n�"C�@_lc�֪��3���3L �G;��L��u��D�ۏ8h�'.������P(�X��(%b�;E�������;�Xϼ��R�S�ZB~������^Fj-�_������v�-�CpAIe����ق�p[;_�D��b�����'�٣��?��-sژJ�l�ֆf�po{Y�%-����*iZ�p�d��e�z�5L�Q3Wk���6�f�z�(T|�wi�ySx�H�����`�мm۝�z��x�r���@u�;��l���g-�?X]��]{lB�����Ì�,�:��A)� �B�4)[��kw�%���ԩN��E=�m,X��.���S�>��yH�c�AZ0��@��~r�ͫ|�����j�����U5�={	�8�;FJ%	�l�=oK�iYR��v(Վ��Ll��s����_�h���RK��ئ��R:�Zp�es�>?�+(�E��S.�pV���QW7���/m��N��I��'-cUs� Q²��F	"1XPq�2,{>�.Y�ˋܭ�?Kub��o�nHh$̭�N]7�B����叒��a��]RPb�V�t�%���@�jv���m^}�{�ǜc�2��ų�Kچ#1��a��������':�s�P	��M��-dq����B������P��o鄐a�4����0�v�$����4XAd�	��E��wI�������`�ʁO��}##��I6v�����*Y��$�^��jXA�q~KM��吝|Ĺd�"������o�O	c_�#���N�='o�ay�)sxջ��ޝ�?�zF�,�ɺ߽��!�~��R(yAO^��	�������E
�H���}i�Í���'^~�T>5��v[o�fj��h꜂<���zO�����>OV�ʇ���s�=�^u�EDx�?¨z����'C��ł; |����.�zO6�|�������n'x�Z�Z@bx�:\�E�*�KV�K�Ϯx���+��4�u��u����{�_,�ܸŦ���7-5��+;B���fTC0���4sƓ�z���c�@���������T-X���H[�PZ~m]�H�Z��cL.��R�\g��6�����YJ��nCM~��.�=\!�O�>fǗpƓ�l�M��N��ꖱ
���U������Z&D�7���Y
�Ch�|�C�*����W5�?o�L���d�s?3O�Ű\/��7T�萭������Uj!yKX�;W���6�4�����[��>2h�����23:���5�8[ 9�xb~g��7#%-�7��K&�5ws�D��8�_x//�2�S���_c���p�����Q�+������o���kX[Ճ��yY�u$��5��ʤ���^�i� �%�rm�C�������!�焎V'/|�4�n��B`J
��a�1zJk�ZFt�����=��?F��&��TbPl��}ke��N�a�~O���}eU��6����nĮ���뇘^Fiϱ���P�T�(�|�c��	+7U�x∉\�(߂�/%���)��{]��Ч��%��2|-��c�P�M"5D|��������^%{��Ɖn�@�S��bY�13|ݙ�ɈW<��v;y��\�4j��3F�v����ْ�� E0�3;�Ca���*�y]�3ey��I�DH������Խ�?��$�B��D���f��OZ��p����oI|0j2B:Jy9+z]��Z�*O��d�z~�O!��1iC~
���hDC��O��v�|4=i(�*5h��@*�Q$Sy����+N[��2t/�֘�{C�Ohn�&͒��"O�(��z�u.á5ǘw7����y�����Q�:��D{��4U���g��������n��ĥ5�+��=7B/9��0�v��kB�d	���o:�Ǩ��p9S�]8_[S4���6�7]ֽb���a��ݚhψ�V��QS�����1+�Wf벺[��^/�Ԣ��x0��U_|��;�H*��{ɣ&�,���>2���;�ǀN;�D�ۼ^k��٭Ln��I[�555�(kIQ�iq�=km�����E�@��h��#pڢ��1�x=�T:�~��z���| �C�+����ũl91񃷦� �$-������W"��[�GI�z��y�P��g��Cp���ցӘb;���oo�j"EOf��~��k��;�Hu9C��T�z��qΐJUL��8�d�z
�{4q���y	 �@�*��h��*�d$�v�mmW'��$��y�)�a����$������S<^A.B�.�������TQb�f��5�Ň�.�x���{�����"�O⤝��-�<�_�[��ADF�� �����hp��SF�l���T�~�ƽ;��(�,?�EƊJ j���?�j.jNCߥϒF�W[�Q�ɀ8���	:�}$�e�-�xq]p!��]�_���yp�z����<|d��e���Nj�?����T>����ul�m���OI���T≡Wl_���ZyIw�QU���pK
����"���h���Nf\�!��jGn���~�6���X���x.L��)Dm��K�'�X�9Y�:�Rg޾a��ӫb(>'�i��.ģ�%.	�L8X��?;	�AM�s	s�*�B>Ã�;�"���������L���zb�*	�@܋Vd��)�"| l{��
����|����ȷ#P\���,jH�6�0���Á�����Bp��Ծ�av�p"3MѿWS���cudz�RX��0C�x*�N����~��f��>;1{�������x΅��@�� ����dȥZ,#X���p����4"/9�@}R�i�x����� ��s�@^�3����y8�Z��?�c`�:�:-"O��2�*Ά�,ԭ�t�����2U���#�c��(n�Ψ�${��E �l||<��")�~��p��]�V��z�MN
-�y�$ ����bH�^��RM%y��)U�|#�F�Ml]Q;���N���+��m�o��-�F%V&O}�2��
P��C��&ţcw��<N�͑��:;��x�wѠ^���z�ᬑ�E�T���@�*]�C\�k ���7˝�j����y�erQ|r��O�c���| ݾk�΂Lp���y�>7�:o�#����En�c���:��'��唘�v d�����x�������v�2�i��ۼ^qY���^t�S�x�Z0VݷdR�WN �6¦�:)p�P42���6�)��P�|�5��K�i��)�<X��u"�g�h���	G�=��Xr�\+���?���|*�5&��pb�q�6fY.���X�W�'&�����!�\�^UN�2
ʊ�1��,�'=��[&p, ��q�ȃ��ʫV�g��u���m
�1ߌu���A�Szd���E���><o&'鑴}�unBG�3��qk���B](d��֕���D�@���`2B�W�A#��k�11/v�E���&1�HH_���&��h�����A�g^��(�e�)(�_?֬��[i-��s�U�B@^���9S���l��F�(5��FS}��a�z�,�����d���P�s�O.(&�/��ET�.�!=E���M���yr��:;�*&��$��J�A�3t���m�%"�h�ȼ��-l�n<wt6>H��^ZU�`��	�va�G�N��-�&��Rʏ���X���7�'�b֗qăs�k��ڐ�t�Tu 
�q9@��V�-��@u{�z��-I9���N�Oy���j��g�a<|��cZPHe�oXcS��O
�nFDd��N	�� �y�z�i��/^e�@\ѲUi�]ѳU��/���x��c��b߷ j�D�ߠ���.����z����y�*ݳ�����2� r����-L|I�T���T|mĊ���>a������M�։�{'��~ط�I$���B�/�;=�I!`�c�c ��,i?��t��C�wF��Ҷ�,����[�ԒS����*\٢�����~=Y���wL��nwC����拒�x�-�P1�T�=�u{B��.pM��n��R7�t�]���4l�&I���Jz]./����K��j�j͠��`nn��qO�A"�R,��1Җ���~����sԠ�!x��*��LA%��7�P�ܠ�qj^]�j��\~:�d��=�>�:�}$�#���9--I��s�AXZ"RPA�:��$*��|"F��}z�ǟ~f5�ҩq��R���,˄�T��dJ#KP���h��+ܟ��65�'
��I!XU��Ƅ
�4�
ᦓo���Gڷ��?P�0Ά�/�љ�$�e?)��,s���xWh�}`p�6k0S�����-�����W�9�L-'�~n���A��w+�4^���B��?CU��qS_=V���#s��$)�K�?��*o���C�s0=�W����y`pu=�S�^�=[¤�Z 0}���G��"�x�˔�rF�o:�P��{�@<�!B%��Ei����qn�'�~¥����m�mEJ�D��ӝ�:^��6M�dwG��xm,D��:#r�[�p��c�F�[�����鰗�>�˸-9���U�l�����K��1����hH��@���p޵%T��vA���t�-��^�U�Y�xEC�����iŦA��*��`� 4nc�����I[��g}D�@	w��.�b��π�M՜�jߊ�:Ɂ0�D]N���r
.�?�D҃ 0���x��*��>2�j�#�Yv�,��w��.m)��~�)�7m��ۉ&\�- Ew�^�\L�Y��1K(~�Vf��h-�k��Nv[�r�~�0a�L?B9uHx};��V��VCe�O�pq��'U7g�n��O`<cO$|>^XUA!�4�2R�v�zc��H,n%��G3��]"�AN�x5b �#Ǩݙ_`o�%/�,��"�1"�;m��>l{��ō�4�^��2X(�(�Ki�1W'X�UO����n��x�Y'E�3���9���&M������d�qm^�G�Z�E�cr\(ؠ��o�r�2{��Jl�h��"a�`0u!������u��ߦ���Cu#��z8v���<	��\n���=0�ь�Xy��������;=kw ��H�'���g�Ō��o{�R���ԇ�Z6I��(d!�yr8�$�$R�b	�Toi��D\��2w�����6Γ"��$���������σ-}iZ�����	'���e����f��
��7�	����D�t�f�j{��
�%:��� ט�-����ؘ�DxX�C���ե�%�?_����E����!�Y����+��Uv�H�\�O�Z��R��5P���4�jY�V-tF���w�ȓR�ܠj����c�VG�].r���S�	�k����0>���_��S�����Qol���k�gb�Q�n*5����D Ӥ�V`x%�����|NЀ��@��]%MZpZ�
߃@�.���`~�L�p���N�E�Q ���Bc���yDvP��83���q�}`'�#Vg5�fm��uW�ĄD�e=,���
�ۓ7�n=��-�G��[:u���������;=,|�����x������K\Mq��0��f��ۢz�2�U��F�|{VW G{T�߂3�����#K2T����g��)�=��n��C�;=7h�P9)R�� l����Ĺ֢Ȯ7��`�yʃ,nnOL��2��<�3�<�0UB� +'y:�v&�%+`���w	p�_D�锦"���Y��nӗ-ד��Z�������c���N��~@�e�[�+WN�T��_APmVd�=$�M�ŏ�
���l�@�K���P��ls�D����F���
y7R�&@�f)#6C��C�z $G���e���%�JˈE���,�d��*FSrP�
�8��m��_$Xw*>B�F	���-Aǘ4�?������O~�c�ɑ�l���r�7��w*q�U��wY��?{:������s�3�!�ÿ�*Q�=�"&	��B���,����#�U:���S�nn7�� ЂN���m�0�#�`���O"�����r�Тϱ�m��s�t��2�e�~T��q��%�����!4��Bn���%`ك6֗>>;v���P~႔���EjްӒ �}�a�8��u�JI�R��E�#A�B�o����z%��{O���2���&1��
��l�m-Ǉ&F`���; 8p�
n,A���p�yQ|9�{=�eE���h�%0���Em��sZt/mH��*�׶i9�$�����G�Z�T% &�`d�OTYfX�<���O�P�jE���|rw�̠�}��q��J��?UlPmI�?~
m��paX�'FJ��Q%�'����'����P��M}�|u�_eM�u2���Mr���l�1���&=��ݳ��Z�0�7+.O�%�f%�y}��x�mL�<�!X6��ʙT��/�ܟ� G�|���W��O ��'�y�r�J��wg5߃,ֆb.����\��Q�����B���j��7ų�����NK4o٪aZb��F�.��ݧ�n_�!,J����D̼S���]"',�t��7�z��:η�4`�S���y 
�& ���'S-��L����q׳k�62tްm�WL�x�E(�|�y���➻١��e���xzo$g�@���{"�5.;3+R��et��!Ө�`j��IbGp�^�U��{{�J�������1An��N4<ѝ�wfH�j��J�g��E����R�����j��<5��̄���������S�R���{X�f�m���B���!0�"�0��%�Hk��"Z��c�c�`��lP$t�HW U� �D{�R��ƹ^E�XY��Q�@��-P�޿��`�t�H:���3�ͫ��j�=Y�ǻ{���ϊ�r�ь7y9��ȥ��/?ZA���6f�!a�=o���>=G�a�{V��a٫�RO��3�Ty��;���Uu�V��u�ނ�V�U�蔵���_���Z+�A���doA+#��NlC	_�:y<o��y��� ����6��Y�֧DPN1,�U��$�v]ƃ'k�E`˪�?֯��g���Q�@���2���\ჴ8�#��=:u�F���>�W��g�Z+�%{r�H)JAK,
F4�OkN��|Rپ�ӊ��ʌ�̗�tC��Aj#��&�\���~�r�f�u������W�Ҵ��)C.�RL�N߭3�����װ��s��.�z�b�n��;*��Wf�{��Y��=�
�~�"���K��������US �.K6d�������������R�C`W#��n�v����v���]~/*j�PfTd�`Pc�s������������ݘE��;�>�9�%�-�,e��cC?���#Mƈ2���,'�"���^��\�g!����0Ԋ�C:��^ڏ���Ě�)��f� �F�h�:���Yp�dT�>�*���PD��	/��������Y	���V�KE��_��E��WK�E�l���ee�$�q �_� ������\c%9#vppj��He�fw5�ps�u^�-˞�C�*=P�h��$&���6=�/��g�ŖL��|�Z<|��8��খnȄ|�DKZE��*�Î.��t��ܯHՁ��YFG|��[���p�`����J�I�t��Q0��� Ĭ��]gD�D.L_�e ڼ��j�ӱ��5&���J��l��*�$RX;n�m
m6J�O���ê<��ij�c�Vk����jK!?x��[&-�,|q�2v��T�8$s�D������hPFu�m�9���pN}դ��;����Yt����&b�3A�af%u��AFc��(��hx��wrs	z�u���&T���'r+�Ӗ�����&b�q)zg�Q7�v��`��Xɤ�;&^�K�[�j���c�1��a�Q��<i͟2����c�H�'���(8���=�{E��[ڱ�U�Zu�ҟ�)��gQ9��b8��j���/��Z�Ƨ�A�C��	�䷽��S�@���n�Sއ�
�a�yec�AU�豵��ϥ���fBfhМ�=P�)�fXwEI�4�̖�R{�1c ��_�"7������_W��*�@<s�4��lx�z�����M ��G$���S�I�(� X\t�,�ڍ��}�dF��R��Q�r_+Ft7�*�vMNh_����c�:�}�tT���Ü�!MJ)ղ	EIe �>�.b<\��w���ڀ�}.�t��Ɉ�V�w�sDU%x}���|�&ʚX6�-1=a����d�U�=�1��V'�pz�"&>D�o�9)zތi�ؿ�qt����#J����u�N�T���&�+z:�)�Ȏd�g�a�qh$т��u� ��:��~�� �$�C �n4��.�k��@��$I7�^q����z�t��x�h���+*叭?�c��E��+�c"�T�.=��÷[��:}	R�=Rݍ��Kl�8ahs��XM�'�����>f�zZ2�W�FO��\��2�����)�Ĭ.�B�=>�4����oaΥ���0_]p�?�n��D���M�G�<��X�3X8�HQ)2OV���!��� ����φ�<��1�n�*щ.�T�ģo�vIh���f�f����۝���*2�K����a7f�c��p��@�������q��Ugv�N����Ghl�x~��[���Ó��?Y�#��5ԕǣ�`�88��^:��x��Фsƨ�bm�!�ٯ>���x�5�m�T���K�{
�B�� �=K�i���Z�5;t����]��*^'d�����H#�* 4T���|����7����Q�g>揾�����#Xϔ������X�.f�?po}�	�Qm���~]�4oQKJjD7�"kY˳_3��_.����:q��G���M-ٮ����@�N;rbtEA��A�{b��marf�������1g��Mq\?�;/�蟄_���{����AP�ܕ�:[5����۵Q�8����[Ѿ��a[�N��gT��&�[���N
����Ec8������T�����>��O����Dp"��z���-��c�AU�'2�ƣ��E�\���%�%�Eu6�1E,�/@��$`"o1=�v�ɻqRM��cEg���z���ZDXL+,,�Qd6�(���;�/�%y',�\P��9I�iOAx����\y�[P�{%�E( �VK�8l[TvE&q���P2��/��H}�Va��3��?��Z�W�>���8|Z�	�̨~���a�l��W��9�E���_��<�����I���3�4���d�5bέ=V�J0p��k>�U��Q��rU��c�X�(AZē�`G�0�b�&�1l�P��lN�<�,^g���1�G�U]t]�D�eT�h;4Y�3��0����C��ۤ!ǿ��2�w��qZ ��f�he�?�# x�bh�c*�\���%�}?|d�����2���c�W0��&�Ҩ�J�Ɂ�#����H;���%��W�qY�ܰ�8���Lܪ7>g���:	wGIk`섧'6qbd���Q��$��i�d�>$o�;!��g����p�����a��u\��&d������2�.��f7�����R�xi�'�8�U��E��6l��ۦu���i���F� �WOhIE{z�b���	M
�����+��H�C^��@z���*�}��A�KW��_=���QO�r��{G���o!q�9)W'|�Q��,�K� ^���m���8_�iڸ����T�A����|�b&��P���A���LԌ�~��f q�:t
��'p��{��e<h�����'�̮F�IJ?S���%�_�$�z�#���.�I
e�]?�5�#��aw������r�2\'Eo�p�y��w�75��R�3(!�ƭ��Ӧ��b+����2@��l���V��Φ��sbA��U����q��I �nʓq��ùt��Nμ&���D �==���	��BhA���!tS�R��5�W�$�#�(����ٵ�1��7U�AJ�qڌ���uդ��4RS��ښ��@��={�0��-��9�%��_�(�O���w�u���P�Wb�,��:����Z���}���ډ��e>��������ܿٮ����AJ�:����'�@�or��7ǯ'a�P"u{�~U؀�c'$���3�����tW!��=�>�y��|������vt�k{��c������z�8\�����"Ƌ�領(�ǜq���䀠�,w��xf{�1�o�m��}�h����mQ���z�ޢ;�$�R��3�oPԥgq
��YS٩��&�J�Ӈ���7�c�<,�Yw�<���&|�O����L�N0N�ul�}Q�`Pv��7�ck j��=�L��W�}��g)�y$�g�d[���=# :�����H��C�_����Q����r���`�s��T$ �g�����JV�_Y������F!���v��3	��Q1b�K����+�݊�v�	0k<
���cr�&W�ly&�>\��+��&�����B�����Cy^�Y�ꗢS�6N����JX�AM휦O��M0��)\����ҷ��-����@zR$���c�p����k`��T��z"����XL[�j}�dtNN�Pg?��E�k���2M���9�aj����)��+zz�>�q��o�EM�~�T�gs�Z���:�*rW��ף�c��3~[���Mk�*�Aj�6��?æŬf_cpv,����`�/Ї�o���/� X\%Ÿ�s�N��W�M6pV�şe�x�_����WIW��e��tNNQ�B�:���U3*.TB�,�/]^z�f��L�����TW&������ʒ��cGU~*s+	�R���Bd�b�cU��e�)���Jvʥ�pؾw��{4��nb5:n���l8.���2�Z�<��F3����X�SX}���J~�!,�ĕ���I�x /Ф�>Qv?6�!��!�P9$r�Fܕࡓ�<�2II9DC����xw�	C�vL�K��%v�hTMv�7�����h��)α��oע-zR�R�*��7b�IJ�t�4�h�^�^��5.�26_[�p#���־��V&i<x
h8��������*P|��i|�o䵹,�H?�E��%���C�aҎ�jS?�����W�*V��/��#9��_%r��h���#�g��[#;�īX�FLm\Yk�<Պ�2j�����&�N���q˩�\c*)˲�kК��(�֡v:���2��3U�˞~��{�d�l�^���	�|����n�"���oZ�o<�>�-ƥ��
qұ���x��J��e��/�F�欮�7(2Ծ�6;�߮�V4����7_&��]�aʡ!����~ζ��1�r�%�d��M��y5/_0���\;"�M�l���}�����S���	���t[x r:d��C�ƴ��(+0��,,h%�s�q`�YR������W���ea�/i��v�!���ʋ�29㒈Y����d��>��e7V(|y��B-s8��@����瘟��
9��.�Nb<2�ڐ���~Հ�C�lH}����㙜�"u
 mB����T��!�x-g�g���{���Q�P0Aq����܋���F��vs ��'7��60kki#���tU����Lj�K�ت����ƙ����3;аtכ���J��sh�r�h3f]i��ƑY���qպn��M�ʠ��l�_�Bn܏�����q�N�L*ŝ��Uq��kBDiVz(*�o�D�B�u��G+()ӓ�2�)���7j�_�m��5}�C&4���qI['�1ݰ{ӛX6ֆ�-�O�k�<'�c2t�Vrܰ#��#�_1h�oD!4��qV�J ����?
Tz͎&��'��]���6�j����zb*Q@�+��I�
�|��B;U��0�J>4���s�����uR��{(�M���w%���_��^	�2��DS+��[g���X�:�׷��D'���3��'#���b��ٻ�"�Ů㞎@���֒%�O}5����i�3<����A\V���c�n%�A�0wQݎ���������MF���D������T|�ej~ L�.�]��S����-���F]n��]e��"G�v�d��8�|��3H6��J\a�$����;�8�Mg��u�ǧ�)�]��kE������I� t]��Fǩ���e�?��I�9]�R��D���!�dF
z d�A�Q�K��~�M�,��&T`�����ZVvum��w���6�hXL���=�m��Se�//a��7b��y�ϥ���V�B��DP��g�C���oUwoX;�"Yr�z>�]7:���R"��у�(0A\h���(5������3���6�M���xa��Ӽ��B�ݹ���/v�+-��4}����v�5����1��Rǒ�Yu��	/C6�_".V"��n�<��hĻ)W�Ж[y �^�MCo�KM1	hE�: +�/u��X�1�w���7,XR-b�eS��4$�dn('M!�"<=m5�[��VPm~-vԣ0�I��f�#��Q>P9 ��xa#� m��&[��J9�Wћ�>��0ǈ^�$ux�L��G���2j���u-��m�/lrr�\6�}kL^fq�\�.D��@��J���VD��}�x�Z���}��0���oH��k���u��εmt2x���m��N��:�����].�E�pK��'���gZ-�F���
��.�en�m��ԛG$�TPjI��oО� (���@8���#��B_`�f9������u���F2q���E�-��K�=��y�]�'�EI�9�!���@�F1R̲��f�s%6?�>#r�XaӍi8��&B�q�OڽS(,����r��O�B��!�A�$t���`V�l��ي�v~)`O�5��t6�Xz�'{��8$��ŝ�7�!�j�miE>_�3��@*ę	�@3��}Դ�'��`�{�]��4�V��]�|
��$y��E{�Ԯ���Gr0��P��쌿I��P{�ӒF�嬝Ʀ���lz���.$
B7����4�Q������/5��E�+���i��(�F���R.-��`I�꣋t��Թ�7c���D`p]��L�I��ڃe&�fO�	��l���pj���fp��P��?o����p`��^�]@�b�5$m�Fh87y��H=Y������ ,�&2^H�H�C}�s�Lc#QfRq�Řkh�?����.fc@�PV夜9���^P�/��?_����2ձ��/$l�G�/BF��� �o���s��㟶����E�~rx�/^��u���-��=�y�@�I��Ű���KKFEq�M�2o7�����Y1-;dʙ�X9�y�vVW�u�%]>����ȁ2e���q��ᓉ���
����&l�xV��R��XI��l��܃9hʌR���I!ΰ�.5���G���H�Ea)n�O ��*!�h�q
;>w�`�L'�[+8w>Y5�II4Z�}#���,`&[S�������z2����5r���*����M�A7���P�,�����EhW�����Q�/1 b�P�x��/�����"g))j
p�A�#p)��q�Ȼd����9 0/~��;�h���T�tr�~�*t�-������ŧ_/��fi�`m�"�/�)0=�:��W%��~� 7��8��-|�~<^�Y�:�54g���M�JP� �*\�0.�d�@�q{������M�􈑤[	M�.����*DK�����Â%>V��Cxj�-hM����OvSwؠ-�n%��\�}���c=�ֵ���";��?F)���(e�VE"��v	O�1���l�qN�-��k&M6?��T �L���ބ�)��&F����e*��|�L������t�o�7�������`��I���g��=K�o�֊�+�ab\y��$H��A�C�y���9SaKt�o��s :Ra��bi�c\ <E��S�nBҽ&2��ⷲK�ߨ�k�&v�10�����Z��䮌0~l�$WZ�1 4Y]Ig/����s֩��&�^ �G�v�>7��K���S����@v�aMb��~{;��ǐ��ݛ̍��X����B��C�%TP'.s���Ɋ���!�&E57�t*)e��=r��D��ߢP������ɴo�v��I�n�cN�:p;�z��KQ5<��l�'2$�ϰ�^��q��CBM�>�7U  m��C��8�U�L��`wBY�R��j+\��mV���_Ĺu|��*�K��)�	b�F�J�:��@�&_��Kp"�!N��9xh��ɫE�w$FFɣIRj9HAr�,�̛S6�=	x6���P(|�b��
|�����+�\���%�N��_�J#Rq16���;�!|~|���7��K�L壮�^�pd�63!Y���{5VGx��1qN|;� 6(�s�W��9��p�*����)��cY��iV�%gn�萭жߏѺ�E����0d#�N�Kq���A��)2�DĽ�K�٦�.�u��z'#(�#��"�^ 1�Z%/B8�����6�J�ĩL��~";�!*���̲��qk���\��H3������RL�W+��T9���?��E�˼�v�(�u�K7o����+%��9��0C���X6�hy�i ɾ��3�i,*�*P��QKz�����
�BN ?oƂo�������A�3}sb�+T��1X&���6�q��0-��-a�90c�K
���Ն�b��O��\�O��D�?iű�Lƃ��1f�����Rj�-����V[$�!��r��fF�&����6��̰y�է��1�JS:��8�̩5)J2�Q+"��0�����j��+0DՇ1��}d;M��=�u*7�';�����mـ��=<QIɝ����a�B�sȉ	O�9{�'@"��kh�������u�>�iS�@.���K;u8�z��s�'̾ �}qB��l�V���H�����8�r� �'O���N������ 8��]�j�[o��8"K�r��[���Q|��*�NƓM�/��3 !P��V�5�8Kl`�����&����Wi-�ݎP�N��?�h�}å�Ii\��0QV��>�
��1Զ�^�:����.u����J���4��mE�C��d�f��կ�����j�+��gZ88��Y�J뢰���j�J�2uR��;*r���%K@��߯U$�F��!Us&�/L���o���(�b�:�uZSw�IPH��A�:�x�3��( b�Z��P٭J�,���|�/{3,Yg�y��**��R�]���P;�㭅,��g�y#q̽Q@��q�ġWWu���֚ВY��2��]�`��j�Q�[���ǎ���b/����&���r���2�z�=e!����d1�i�B#��B.<* )�z�7q4���aM�ۊ��p���i����������e)W�j�\����U��^�1�C����A�v˒3[�$�Gj{�������[_�oRX�-�Vx֙�|c��pω�O�G�0�(��6�����8� �T1j�<P��̓:7�w�I���!݁�	@�=v��4������E�╩4�86��6��Ct�`�tX�@��%���(�rQF(@��0���ֽ���8C�q-���^3w����'���2����Ҍzt���l�Oc���4ܽ}���C���������v�|>�?��rڧ��t��'*nh�[٪�"�������^s����BR�D����cQE����fұ��H�YD��86�ْ�q���<���� @�/�����������&��ȓ`��N�ۯ��pWrL�ӭ���3z� ^u�x<]6����,^?Bp���VAiP�؋ng<�f|���څyII4tDV��Q�J�,z��Y��}�B"� RU����\��7�Q#�X��� �*�ɕq�s�+{�����!������ ��Z�$��P6]?ÈBwN�_���f�Mz���!�'(z�*O�O/�A��h_��U�erY@�O�h�^��gk���<W��:>xP*��!�#k�������fڦ���D��ќM��F�8�e�<��q��JX�Ir�(�.�����5'�Z�)_�a�<�,�I\h,�����Er���f���x�=�7R���@�R��C�1�
 �P�y���7�	j� GO����}�׻L��7��m�x���n�q�p_r�4k�oپ�*"J Z%X���"���R�8�����%|���x���k�Jᚲ,8.s�A�=
'��n
m������؁��hnGh�tr�����z���)��3J��E_�W�Kz���d�S�n=
lb)��8,a���.B��wz��޾u엢6��(�>�/;��F�JAq��e���%��3�k�{xI��?�y���K��m~Z��[���*�tȵeV���?P����n�}�1��]�d��Y�4���VZ-��LQ���l=o�7BI������D��_X�t"�`�͚Zf�+��J��g�T#(�YT�ۤ��� �N�y)���W6P�s,)���E����
��F[^*�'���.`r��g$Ĕ�c
�ܪEL�}�Ei]�T�+�д��������'�'=�cN��=`]P�|��X:�J��`DȐ��C�+ƣrº���R�eY��E���B�Sv�r��D)Sd��tN���j(l�[f��!��X���h��6GL�-�XA�u[ʒ�ćk� _�p$}��eɭB�^�"�怜����N�;�O��*&ו|ʞ���v�[נ�3��1*!!�G��Y�vo�!@[�GX ֧Q(��K��"���ʆIVO�����={�mx��u�,N"b�����l��7�����6D�Ч"=�T�|�$�� ������z���^�F�m%��Iy���9�����	cu���Ә~�``�ƵւV�X���*]���o��+ �+A��o]`&�d��9(fg��`��8��vaGDyf�K��T�B�(>R\��y�čw�����r��ۈ��ȡ�w������%��1
���χ�9�nyܗ�Wgx���]��%c�lH��)��@������g2�c�9u&@메�3�T{{�#M,(�=�d:�ƅ#K=�����tp��HQ��^6>]x�뀾��8-����i��9�cB43<��8� 	^�t`��@�)5�rae��!?zƣ�>����e�
��{$�"{���ԡ��̸�<�Qx��k��^-�z������Li�5I��������q�^���ג��MZi,��)�������mn�w�#�s��M
V�^5��4};1��}�'{q�5�j�ttE��fVp���P��>3�]�c�=�w�U���ʾ�o�Z��v���w� ���p̍�b̔c&
�|�� �O�u-��VB.�ݬ�,�d�Mro���7���˔ xD�W��'Dī'��49m�	1��@�u�q�J�`��!u� �C7�X9C.7֩��U֍�m9�3cD�9MЙ����������<��w�rGGVՋ@�э@;�Ψ��h�i���d�W8[��r�[|��{�	��M�嘋ޏG���mĐ���x�OJ2��w�Z|��s���fZǱ��](Ĵ�iy��`�ӑw8���oK�����R�W-L$,�n������ን+95�fjО�R� ��{ݝ�s$��O�ټ)X.�Y4������.y�����T���0E�U�Kj��0�a�2�0^	�p\ǈ�RW��A#���/���cl�:�*�����]�s@�]#	���fE�Q+U
��&���)�#z�F���wT"G�0)��_!pdM%;��� ���6����S�Q�Zo�����vg�N^�m>�j�0����U�{e���ɸ������͈'�H���\q��|��sV�(��7�v�U��q4c�C][#��d�p�M(�P�<���{5�� ]l�*P �\Cq�LN��.2��g�9&xf
�Ʌ'w�2��f�{0
��j�U�����4m�����6f�%썥��� %��M(�֚,�9�؛�!{H��c=h��Ka�n�[�_�ë�*B��o9\�d~�䋲Z��z]a^+����l�q�긁0㦴�7M���Ͽ��Q���e�lʀd�T�s!�1U�ƀ�ڙ���%�`�S��E��r��rm��lPP>=3����T��mZ�h����+�˧>�{8&G])͡�*Q()N<".� ��D}�;$'����D��M�f�@����):߾�������HO�,i�[��U�a��ԯC��_Qo���پUY��tNv��w�^O6�������������s��g���:V���2=��Y=ױ�@c�K�G����V~��?�uKI9��ij3�I�;�KV�8\8�da�6x�_�*55�(,�)�`����6�Ue�ю�de��lI9�l���F깙E�MY�����DH>fl� y�v^a����1Y-�D���c˒��S\�in~ck��Y�&��6S��Q������xM���f�D*�Ua�� ��X��Jj�\DY ��mͲ���)3��P��'�-��ţ��HEFe{�H �����[��0��pU�+0�؈D�o���7G���⣾đn��<Ǌ-G��e�	��o�x/�]�,���Z�#��0ޢ�*��/�����n�]�1����A�7�k��U�v4s®I�P���=�^Q	[��1�MǠ;�A٨�#�	��W�� �����V��Z4>uM���R��y�	RyE�C����G�h�aQ`Ks\|8�̴�+���l��cK�12���1ܔ��C�l��7D�TW �Ď�?[�b��c���%�v�v8�{u�E�[;I ����{<|
~2M�R����1q���TKv�]#���Fy餂�~��W\�@��G
,@���b�k��t;�_F����ə|�&��ƅ�h,Oa�Ϙ�Nrh�d��<=Y~�:|[~�}�l�C�I�6'ȣ<�������1o����]"��
�`\E  0���b����J���XH��8�8�����Y���D��I�X���h܏Ԟ�]�^�o&l�6��B��o�=Ig8�8D��q��?��nwp{3�]`��h���}nH��҅3Z���e�ȟ�����5}lo>�9�����`'��� �?*CzAb+y������0</Fp�y��#d�lm ��?=��i�nf��,��$_A;�ކ���h���*<|��Iy���[i<ː���v��\OoS?�[ז�r���X,�Wl�����^AYI<��t��Ym��-�Ȯ1���S����b�行6����Ñ��d��F(�|�'6�I���ɬߟ����#� G'��l3e�ۇ�&�����U���HB���X���nj����#X��,���)�/����Y��nh|h��S�ψW�0���Z<-��l�#� ��鸘"��i&k��9"kk	,����E4ѱ;�\�4��X�*C{���m�8[閟�靱v�2����3T�WR���'#S��h��د��.��<�#Ɣ.�{2[�g�YŘǕ@��-Wń[�4a�=Ez��ʖL���V6�٪.�.WY¡��h�(,�8v��gw_��.���x��I	�3XO����M�Q��iA��1��	�ق�1܊i���쫵�&H��s6ϳ
x>��W|ؘ�	K3N�ZZ�L�l>����H��&iX��5&�58k{˅����Њ��])���lTdC�~��8�%����Ax��"h̭��Y ���p�����G�K�����aF�P�|WP�����|�r:&���AL�n۽�/�g�����u�YoB����
���`�6��g��<��x�� �!n��^�<��)�31�������Mg!:f�mJ�<[k�%X��5��0@�D�j'�������s/�|�X�z��óV��䉃X�ɿ���p���EB��E�%mepN� L4�eco>�1�˚�d]�5Yc�ۮ'L%�0k�s�����{JG�H�z�M�G��&m�tn�W̤��ơxɹ+j~��ՠ�$� ꡶�aY�Tܶ4нgG��8�.�+�����n/�3 Hb���.�[�%�U�#=�q/u1����� ��d��~r��E��H!�&��X��'c�#���p3���A�N�ܙ�Y��Oi���H%���J7
 ��`sit�A�sO������#Xl��}��Vy��2�Ip�ȳ��v JNc���N��5�6���Сiü|^���C�7��yp�P������&�~����~lS��VU�ׁ9�N��^�I#�l��[�ٗ���𜢛I��o��Ē��u�:���P��L�{�2Q��i�^Τ�$
� n.����S�ٱi��KNا��`��SA�%:L,�����d��ּ��[�(TZy���yQ!B/x\�Mdb�a�a{Q����A8�%8��%�˓��lyeeF]�[���c`]��"�Uv��}pn������E|v�$�������z�ٹ�k�]:��u�> ��U`~6��*��F>Qh�~0�,�+����!�=��Y=��$T��{�8X�,w����ޠ�X?��>8���)J}N"��������#]�����&��G �N��i�,�0U��A�F����8�J������̍������[���%���y;�i�F�U��9��y�JL-���1&������ϡ�,�-�v�,q߁LoQ��q�-�ża�N����AGĝ.�{~Ϸ����".o�O�a�]%/[��.�a<`̻uIZ
G�ҥ��P��S:^�>ADˣw;g�FR6�T�2],��ց`\�V�����C}1���^m_�{#��'@�5p++l��Ǭ�@Ÿ����d"M*��3�\�=^xh=����\�Z�� a�,ve΍������1�y��ȵ憨���|�vL��n�̆*Cn�s�S�7�N����ܠ�6O
(A��R�Y����-�%��@LGNi�R���&[i��+�vN1?)}�q����9�~� ���Y����2����G���1+<���jy;��9HS �:�&܁G��H�u��;7PK���9�+�q����-G:a�9�#��F#2�A���6�f)	��V�_�F��$�~�!8J	�� �K�Iu�����h�VQ�4�����n	C���A�o_3�{i�ZL�Q�㞧6����3m�����kH`�Bc���'��*��8�ꎉ)>��,2c�d�gȖC��F�>}��kA�z�7�pȟ����2*��?	`'�)MTtD�[�^ã�ͅћ�F�'!7��)�}獰��������i���Z]��P�2�	�T�òQ�Xr)
�+�,/"��LGWwNۘ� ���<� �� �����������͗S�=�u��#���v�F���܏�-�͟��/���<K�&���*T�c�"�5��k��}��[���8�^�?�E09s����_X��flDAO�ܶ$l"�HN�9�YV�d���9�PB��Rtd�p�¨�c�<2:&>��Y����/�}eN�3�VB�7��A7�t�&	CP�Ɩ
�1�8�#`� �����p*�-����=Y\Hc�9�K�`�ZK��J^�MՇ��v�gB(���v~�a�
*�v��&���U� �+�����,&�G�W���G0N��F/���貴�^�;\0o�k�e"�_�~Xf�)]j��yw�2���w�`�� j(����Pi3	D��+���+����J�1�$�C_�?�gR�n�$}TS'ݘ�d�+��No%1j�0��S�2��/�?NB� �p�I$C�=6���w�ern/
������e��b�������+{�?�~ÃL㎿'ɓ/�;0�Y�:.
w��[P�Y<�b54ܠ�_�E(d۸��C���]�-g��`����iB-Y	5	Q�&*n�:�iA��?1�"����xY#���Q��Z�$f�}���Q�ܛ?���l��#>�	���e)��8�8�f��hQ�٪�/!�^b�nוa_���!�l{X�%�E��5�9���q�U?:~&t��Eͮ�H���q�Gݱ��̼Jo�ϡ�7���'  =��D�
,���dȼ�k�}�3��Y��dA�ۑU��-WO1�l����C�p�8k���0��uD��e\�S��@�A�PY�}�m�I����Z���tbaq�,I���t49���{�O����j"%�UKLA�E����械�Y��H�����(��`"�z��=�,��Ķ4���g��	�����p����9��ޚ�N�%э���rJ�ڪ����ݔz�D���`�4�b\��	5��E���R�H�+^l�ꆢ��ƾ��%����h���U�G����M9>�xrq�\�y��$��̹݂[sZ�Yٙ�|+�y�!�,Lh�l~��}�E*� h&�:`��;�ɻ���A�(�Ç���}�-�+�~��TRkΟ��n\��mK:/cj�p�)X�F/+��X��T��,����.����Yo���0�_j� �`���T�
��ݧk!l8��i�Q-R��U���}<�{I�-��N����b�Z{1$���4Ŵ3�D��P�D�/�'�a̭n�4�u��Y&vCe�@؟oM6"�nT%��~�G���8
��q˰=��V��C~t׆P�J��+41��K1;�]P�v�NX�T�E5����X7�G���wA�ɴ�殺�Mͨ���8��pɛ�Jh�(y��ߥ��籴J�Ʌ�yɬ�}`:T'A�Hh*�3����y]�Kc3���1\H3X�� ��U�݂N���`����>_a��7���d�Mp�`,ADnWLd�@��G�wA�t��K�{!9%��{zy�0�j�/f�n�w�g��_5��xއ�L$	��	՗D=�G�^����n�E��i:/ea�ceș��hZC���c���ҹE����D<r@�S��;}+zKG��7=!H��c͐k���H���^�u?q��DQᖆ�v�B�wE�k0�F.��}}��f�.%��h�_��̞����2�)B�M������:��߄��],�>��/y�z��2b�2�R\����g3�#�J~�S��A"�03�ꖉw�<x�<�{U�JYP&䎋.���q������D���n��<�2�Y{���7�: U������U�M�B&̋���,Kc<z���u� ��U�a��ŧgx%7�H�S@�u�$�=C�zjd
%$�n��ݒ�|��S��׵�4{�A6����λ��q�y�;g��Tut3��M�r���|�,9^o�0ƪ���L�]���!�X�"ےa}1*��=�� :�z��� T����e���&����
n�*q�O���n&F�p����K_l��Ym5��0'�[Y����x�0�p�"P���h�O�=X�9��ў��8��A�#�gϡ<nU�ͥ�
��пK�c.k̘+�DN��!i���"z�R#��ާ,�&�	.J�Ó�#R�\�'����^GL�"K�n.�����I�P�yEH&��D@	��%�l7t	�2�n&(*?��vJnȋ���^���nG�S�ح0��8v����m�̿�K�*�ӎ�z�Ί�a�e���?�RH�+w��J`�|4�i��j�kG@����}����Y6Po�^2e>�1l�[rp�~��Z"�}���!�Q�R��zI�rϷ��K�o+q�R��m��pA��+e�S��n��2ibֽ^����@�w���!�11�t��$L�4 �  � �T���:lj������??%��� Yi�]�9c[�zp}��Md�M݌oZ���M]����(*1  D��$�����S���Y�~�Ŋ�Q��f�A�a�!W���QodC7~�Hh��j
�D���@Q&��o�rR�j a(�w.�����s�I���C�)���m,.�6�[���a �=3b����m@�����)4��O:柭?�_�0�~��� 	k�W�ZG�7�d?����p������<:J&PNΛ��	�xuu:�#1r�_t܆V�iQ���C��*�������8,��<!���*�D�8�m�ڸPP���nx[��'b�w~β�V��<���R;�?R������7�(��`� 'q��t9m�Pp̽���n����&�����_p�)�~�/)��N?F�WS�����ʵ� �c�_%�>��>��I�ߐ�G�16Է1|�S@�#���''��+��a�$p�����'�4��1ڄd�t��~��g:W��h��]nX�,d��h!nZ��f�E�J�&
?��6�0�zc�?�:(�3+NlL' ?F�!7qB!��&�	�5��k�� �i�ߔ���ԥ��ep>s��Q�w�7��P���__Pk��Β�C< ��F/f(CI������E�Z�K�-�_QhX�~.x���i��;�XJ���s�`�p���h9d��!��qWMX]>)T����H��L�/c���϶Ŏ�4-�<��_h�:�Dа�:o�k��¨�7B����E5�tW]�C� D�J�W���]ט�i���T�Ѩ��'��5U]�����e��xy�5�Md�lm��U�q=�!�F~|��E�o>�Ml#��aZ�;�?iS�11�Y$:;��GU8��h��lݷv�A������^��U�������j�"t�gpTc��悛�8�"N[�hx��+юIR�S4�}\�S#���D0
Y/5j�o��h7)M�~���Ϗ�%��}�I,���Q!��ER�4Ed��_2�Eޟ8OB9W��u���*�S��׿��Nv�Є/�}�!>�F-�<K�I;.�:�
�@-��֘W�YG5��K����
of��I�
y����Jw�k�A�V����{��)�I�Ƨm�e������W �9L{ó��Ꮦ�5�ƀl�t���HmT�rs�Ŗ꬛K
���t��1�֘)��?�*No��s��^�F�!]��e+ּj�n;���(2	!)��kP-D�o�P�� /��uh�����\PZ��i�������t��Í�>�'q���֊
��:߭��I�aoI���z��L���Z��f���3f��-�����S�频�"Uy�E���Lf3T�pX<1N�PK�SN��q�� �+����s9�yj�_�|\j�����L<h*S�:iU$]p	�p}��{�)��~��	D��5q�֯b��(����ܾ1��㐜d(�N8����Z$Ww��pȣ鰐�P
���u�w`�{���d�וdt_CA�c�'BO��Ӡ�=ǳy.�X�����*
v�Ol���o��#z�g��o]Y=��"��M�9��y�/֑��$jZ�jN|m*���k����!Q��3sAY���طg�%��:c�)?ܱ��H��0eu/^l|��Q�o���}׫������,6]������l쎋��%�I�?q?y�j�e�U�g�:v_q���]��ȉXO����_�H�ᴚ��f[���?*hUR���r���"�k���I�k4)���)(�rj�z/�^����O~F�Ub7�ɂ�-�X~y�Uxz�c9��>떃e��:�~VP:�S����}�-v�tF��d8�X�(eH8����wuƪ?���ːd1>9�LK�E��$��xM|4%�Bʴ�b'5,<�	���A*�}�j9(w���d�-�<�9��gez;�eIR����|nBOY?�VK_�~�b<l�t�OA�Z[�V�iSI��LJ��āG1DD��;9d�E��?O�X�b�����Q����ɐ�5cpn�]~�-J6�c�9g)Ny�=��� ��~P,�3����+����3��g���}
rϫ�ad�(���J�9�h�� ��A�:=��騈/c��)s*�@�Ђ�{x�������	�fn���%
�@s���e�u��zKŋ�N�^��D�q��'x�M�a��/��5�ǖ���+�0/��`���n� !��=e���߹أ�x�/3�D�|�p�Q��{�\�!6���0�s/����9�=���R�0��� Q�>P�+����]V�7��//�fw��1:����P^G������WZ�.`W޾��g�+�1m��8�����p�]��MG�os<������w��g�(]X:�րL-Sq��	S6��P��T���ǇV��,��4-_!������8��CR~&�BŠ��	a��]���XG����6X���R����mvo�	�B.cr<3�Q++II/�O2�����g���f�_S�>�v��V�1�H���Y��jH0����~%�i�Z��F)z�_���+�Y���jQ�eb쟅Vc��V��/s�b��Y���������`���q��l�+��yv*����ax��鶹C��,�`��^�����f��6O�\�6���}���~����χ�J���fq���u�y��<��7z����
￥1C'1w�����::������9K����F(