��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*~�)���>w�f�Su����cϑt�ڪ�,t4�EЖ�u�Sߒ�ޖ����,�ĩ�M$0"�R�~0�!,k���<�]H.I���"w�Ȳ�(�f	:&Ca� ct`�Qi��v�*�By���Y�9��c@&-�GQؠ����SA�ɐ����:jSKR�D,���r������$鶴�����X�1�Բ��I�f�pE�'M3T=ю���_��]�OͯCf����^�E_�
��t��/���p=�qz��?�@�~N�;0r��>b��Fz��U=���9��8s���
=z��w��k��4^��`ߛm����gt���S��.G�=�[��.�:��<B�J4�soM,��}��b�N����PA���<ԁt�@��	�a;���inN)A6���&Z��c>M�&OS�1!�A��y`��X<����&�JP��kS%=<�#�KRK��(Q��>Hӈp����֩_k6�G"����sm�X%NV�}1�F����L�r)���ǜ��"�j�v�����5ҸN/�p
��� :���&��&d��^� �X�GG�x�et�Ff]>jA�>���h�a���KT�16E}��`�i��J�k1���e�9U'��(�L��_�X|y�J"�j��f����~"u{���طP�S���QY�ua�u6��8�>��ఐ����b5#f 6�2�<D�E�3�T� ��Y� �'�܄M�c��q�M:Sgt���j�)�#�#��d�Y40�ﶼ�����hlS�)��J�Y������ k4+"�r�$, ����ނ��/\*�,ӗ*�����^.r���xV��6FA��YxoB�b�Jқ�/0���SC��w��Q����:Kt:�-/=p�UfyJu�6�-U*�Ɓ�uǎĪ�CZ:�l�t�G�~�9�� ��)�qN����7�	7��0����̤zU���lI�`�����h�p^0Z��ME�PȨ�gX�z� Qi�B����@#@>~�>>�C�f�9V ~�CPG��^��ݝ�
U��f��P9	�ÈTˑ�N�%�+��a:�X:v+���4���[�v�bKDjf�pg����sTe����x(�`�L;NqK�p�����ҍ8˕u��4oB����O̟�B� ���v��>���4E�S܁�N�i*�S�B����V�����m:@��e�,� �Xx�N� �s����z�\�G쥴�<�!M:Z��2e��>2���g\����+��z={�]b�0���sNC'M=�3q2�s�%���b��v�桦]>�F��L�*��fX?�2|w��s�6�Ep�7�=X��m��9IQ�Ԍ���"IX��=���#��J�l�����S{u�"�\Kڮ܍�,8�$p��bx��6cO󁸟��!�z���I�"��O'0lal�8RR 8pƩF�Sr�IE?\�нeG[���gH$gY�c��"i5��L�^���\	�W~�V����@��(��0W�b(�ʧ��uO�+?�Q=����niyjs�У�+�"ߊX��bN����[e������+��+ޠm���b+l�8�9����.������n'��q}C�b��4�F�n�M��
���'\mc$r�6�=��E#�y�2�;���F(jN7?\m�?�QQUe6����S>�i$�nI[�+,�����˃�ö������d����K�F�)�t֛?�8{<yOw��|����8��ԅ�^fz\D����ۍc[��pY�f�+͑����̕h�Q7�D�V��ft��b��ڑ	�`Z#��V�}?R�,#���rr�pH3��&�VO�|.6-NF�\�'��tl\G^`����30��`�HW����ڭG�~�r��5�i�W���@�x̎���%�X�¼c��t�f��9Yx�f�bL0��c�O�8�!qBq���u���\��G(��;=ݓ� �B����#{k�Ժ�I�$�&U��ܰ$B��,����R�+��-����Ł�V���~�����+�
p�Ӥ3"�WG��~��/X���h��&6Z���٦D�����4Eb�fT�K�uO�3�j�����i*�#�}8<<Ǖ6@��:�e��ë_�����^�)x:�ٮ�}��gB?~K6W= �?&��^�x�+�oI�r&VG�ׂ4טة��%n����m���R�K�7�|��F����s;��1Z�0@���.#|��+�Q��}(R*�ۯ2�|������*w"��3��6c����=uu���lQX�4.���Mmw9��B��}&�h���'�Fb��\gΒ��S����C���Kb�%_5��V[DXG��X8���<B�N�j�vq�#'ՕkϤ�h�8�F��d��$a�����m��o�UW�A��BO���oi�t�R9D>H��p�(Ί�fT?�{��&�;M_�G�Oj/��a�CS����_d�j�j(K[l$� � !�p��!�U`*���l)���cz��o�$k&a��{ë^5���q�YT�R4���n�Du�ɱ�쐕�#����+M�$�?��R��^]м䴣�<?�[.z'=�Y����J�O��1���Z���;Y<�m�蔭ߢ7TBb�/'�+e�zjh^Xg�G"���z2Bf�FQ�rc���J�)N"�5�ĸ��P�R�_���#�۸���͟Ix��B��n~��� �(<�Ow	iճ}�!�u�;��X�Sz����v�A�p�kԇ�<T�"�a*tw�#h���<���Gd��E^�r��v5oPҗ��}�|t�Ө,x̰���2�I�Ki�v��Ɖڴ�\<��u|��Z���\�I���Cٮ -@��S��c/}�i�t���?�q���L��������c�;�[�~�m�O_ۏ+�mD��UN�=��q� ����@Á���wr:��PT�X���d
�������#�u�h���GD,�G�xĠ��� ��V����3}�;���*��옼��,�"?|,�F���w��`a�k�5|�:��k�� ;�.H����K�s~� Hm� �֮9��]�pP�FF���MWU����� �w;1��d{�zk�&��Sb�I��i��"֜$g"�b�Zm��v��D�j�d�
mT�3��C�:�r�j*֘L�^��x�kܔu3)^⚔��p��l�?�y2��.����=�ҾΘ�f�aƮFU�LO�䂙[��*N��7i15k�o���H�" P��R��BhB	0G��}q5�tӄ�� .�b��Vi3�v����낞p��#���b�׋v���T0��T,�L����e����q7�`�7�6Ɂ��.�l�V��Uhp�h$b)nЮ1�ER5?�{k��?$��*-�����35�7���a�t�!�A{�<��+��_�B�����֋3�D���% }�>��Z��^��\���/�Ø�j�V����<�	o�-�1EHH]9���Ut�e%(".������9c�]%�����-�/��������u�u�W)�����*� `-6M'�"s����]�(�p��8�����X���϶1BU2�����?����T�{�Y.<7~�
�H���TV_�@'㩢
Ri�� ��h$���?��h�*���$��DD�_�k��Ϝ#c�4����CS���)��o��	5�h�4���7��$���wt�)d�����3NN+
T��f�BE���$���)y 8oٛ�c����f��:\�����7.��V��L���p��^H䌈�Y��5� y� ���0�nV�����J���W0f�����~ܳ�.,k'�V�� L�T�؛/��'A�UF�4�Qڢ=J�h�pY�z�Z�A�V��\�M�jɓ �6�8�������bF�Zؘ���w����I�Cc�'j�U@�<�P��#�p�q��ql��
<p��-"8�H�ğ�DȠ��E���Hȸ�,��0p� `.z>2�A���+�-��n^���vGT[
F��i��kK�_��Kr912r��o�N����F�e��Y�{��l�82gf���7I��?�.������r��1��������Z�{��=~Ptb?�#��[���9>�)��&g%䖖��$�HO*:u{n���)^��퉿���������c���je10�ԋ�R�{0��O�{��s�ʤ>su>s	��.�7�|[0�ؐ=p����q/�V Z����^��r��%�
��7y��`%�Y�m�W���[K#�9�m�#�Q�C3�bu:u�|U �!�)Oa�9�O]���5?>y(Q�����%S�m�Ǩ�~"dF����Ӟg۵��m��Q(�da�J���ͩ��@�
۠���-FM4I%�����hIh��>#� T��+����+^�\�htR��/�hn	m�,&V�����"�o�50qh1%��X`/��DR����IAm"3%b
���ݦe6t9-G�t#�ؐ��P�iʃ
%޴�B���}�+��~eY�u��Zd�Q7���,i:;��K��#@	�&�CD�MH�r�ZG�g��-ŗ�"��� �r�\<���
�L�y'���y
cf��a�u�X�m�������Ǟ+�N� ��p��<L�/I(��u�-�D��8;Ȁ5/]�������<��K�64��Sf=(_\ Ƀ��U5c~��4z-N*��%��!��&pU�IE�N2���g~je��w�h��#S������S�U�}ϻy�z	{���ԁ�]@�s��i7$v��xw1��!����+ ��.��]"��n�æ��İ\|D#���(_�K^��O�Sh8i�e.�z�?^h��B�7�Q�I�E@�ʘfLE�AP�8�����y��M�����	7�Y��ޥ�S���w�R�"�y�T�:e~4��� =o� }�}�U���|OU��Z\?�,9�2��J�OGYzYf�'�V���a��3?e�@VG&|u8O8��R�r�u$��G�[|� �ܥ�΁�z� �X���������2Q�hl̶:0p�.%��[IF�N�W#T�3��FNϡ����ҹ=��+`v��b#`��S ����^q��m���'L�Υ��2���o1�w�V�䘂�J}��\�P�ѼLR＜ٓ	�:� �DC�VVӯ����
��`��^�C3���E��y�TF��7�:=x��Ze���BF㭚�|��i>��:8��#���]m+$��~͜"���$�pTc���2�����fi��v{�_;D=�Ļb�����)�]���u�qi~?@'w?N8�GW��,\V�ĒOGt�u$)�!?3���7Dk�3[}�#��Z�m#��dV[v����4R �w}�F���F�Y\�K�S��;�8̨@����2X	�
4������78H���V���A�)5 �4V�0���|��J�eN�*״�W�/�}�G4�u,Њ�A;t&3�|J�?����	�a%�63J0LD�o�u���rՅXg���;�GӮ�*�'�w����b:��0�Lw�͘��c:x����҃�h� ���AخDC��f&��Ε�gD��":���o�9ۑ��[� aX��m����Oż����]!Q$�)��壽e��s�J�X^���		زWj��[��0�H�Jt耠_Q֫���1���/%��0�""�Y��K��5!�_QW����~���u.[å�X��ιo���ҬCv�!�1H�؅^L��iY�Li�b(1����R�C��q�g�<�_�$m�[�w��Z�c��gP&���S��~�LX<:�#�s�;q���TgxR'Z�0�"V����H��n�s�K-���ҝ��>�]�Y��Ml�5W�������"hjy��~+Y��g5d�h4��B������I'�mvf�8�lʆ+��x�A-K���3�oT@-�#��a~�=�����_3#Ȅyk������+�?0��N�>�?��0S�N����4a��f`<T:��Ү� i���6�����)�*�hN�{m���)�.�_9�\���[ش��i�ʄ��Eӂ+5����.c�!a<uH;�1b�L�{�K�G���ʱh�)��4L� �`[� ��«�Ɩ5��s}�w��e�"�<�Щ�r����%��%]7�S�����j*����f4�ǀ��fTYNJ�2��]v� *�	j�k|Xt�-��I�;={���'F�SS��$�P�l�����
��b;F���R=y��yi��j�T�;N��CK�V��8vZ��)^�h��}���i�KӅ�&�(��.n9�,W��_���s��ܗ{<FobF�+�F�d1�[�e���
6�R$*�Md9���b�Xn��'��v	ڰ	�C\4�RT	R�FQQ����j@�98ǽ;~!j+��J���UGs�Ce��̥���ftЊ�W��+�8�՞� �'Ǯ)���أv �&��cck!n8[\�ǤV����(��K��^�$$�����E�i��Z9Ӏ���;�?<bp[J_��Q���_�8ݹI-�9KWT����&E�w),���'m�Y^��\q�Q�Z��)	�uKz���iZdg/�-���C�Vt
&5�	����d��H��8݊,��E� <��(�ggt2�`�_��;
>�O�Uva7PXhn~'z�{��h�y�����L'G*���(��{�xJ�P������nAx�}���'�����槛_͟j�/�E�/2��Ђ�W&&�c��!p��v^�o�Ȟ�!Es0d-��$���:�@AR*Bs�Qb(����&«�9+g��塔B׉w�	��)w7+�a���)d�R� �ƓOV:S� Uf(��B�P�4�Ӛ^�O���]�S��	wq��>m�����g�>w�ǻ�mjhG�⯤U�Q�\]�ܴJ2yډ�\	����֘���6��V2�&iK�ux�}�~[���wNiCw�\��q|��]������"����n���\s��HRߦ�fŨ��@�<����K�(
���e�i�p!�Y�/�F�i�P���
�J���Ҋ���;��ʤ���6P��=��4.6Rd��.�o 2���[N�p�-%���p5N���	��_<�o��Kj�3$(啗�T�<����l�����tл����.Tz��"k;{��_G#Ivd��E��['b~�������N]�a��U�jf���m����^&��
{�[�$Ku梸��=�j���qY B�)P9����1��L>��W?�YݘB����%��^|��7�y�]ޓ�*^
Y/������Bu��&�=���
m�Y�	���s�5xZ]�@*,�и����7�r�}�ԩ1�+)�y�]������:�?{�11n^�=O*'S�۪�n��>��V����ā	gN�ol_�>p��{@_lu}2p���(C�]�a��%Z