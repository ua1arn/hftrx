��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*j��d٫_u�>�ȍ����"�+�"�sL�ĶX�r�
>{X�oQ;e.2�ζ<F�HV�5�D�Ms.ٶ�(�*��?��$ck�o��Dk�g|Z�Ԛ���S�3���Htǚ��;a 9������;�1�� �a^��6T�����?U�`��(�
c��$4a���IR���wTR��ȗ��� J(b"�[�ᦛ<��!�E��b׵�dP]�� � ��A�jj�@)^"9��@��|hS\Z�@���*����g�XUYlwDݙ	�W�L���3� ����L��'c�G��X��ggl��ע���1��Eي��0��Ƞѻ;t`Ej�����G��yf��¼1Η������!��\������C��?l��u�.���ޏ�*Q�J,���]H?;~'��{]�j�:}�^�i���L���E��:/��]�ߚ,mN=�ys�!�N<qd��?���ųg��
�X�E���kx�6�y�~χ�:�Q���c(!	��C�&)r��^�ɕ���ŧB��[U3q�7bCu���}��Jq�[��=��0�S3l�ۡՐ��A�]d�'A� *��3�����5W�"���Vh�'���x�6w���>Z���q� ����V�oSk��j|Q
r����3_a�ۨw��o�
���� ���Q�dT�O>= %�bs�ᶠ�h3�B�V�ҿ
E�"Q[]��c��M_�mk/����@�j^�
Z�M�?�
�|�t-*CW��C��EN1�A}S���R�>3AO*�2�`v��{��IPr ��?v� JR-�58pgވ}W��͒;Ǡ(�L�%�K�������T��C����!�I�0�:��SY�J�sc��Q�c?X ]K�5��ߓFIz�%�b��a���toE����\;��s8�U$�_����Wp����d��R�e�ׯH��7>�L�C�BR����^$�D��@�$b-	0`�	z����$
Lí���1U_T���}ͅ� �y�_� ��GWE�Y��r��h�`7�u�?FH��b��q���La��A/�M�V Ry���#lwՑ�b�Y(��j�6�K����V�[��̻ ʉ�%��%�������E�t$���BA���{N�?M@�`�h�Q�g�\��<^��
M8�uG:1�~W'�� ���;e��H]�w�!�iQ���3U�*�>[����w=Y.I�4꟧-|n��������_wY���<�i���3<uqR����g��H(��2�����6+,)SV,(J�Q���7�L1a��������Xa��	6�s��X �iϝ��a׮4-��~��WoG�)�F��ίHݶ3�"J"6e��������a/��mn��Q��E��z@��c�Ɓ˸j��m��)��;A?��z��ҵ���3ޟ
��<��T	o�N��5-�W��~CB�X��C'�af ��a�v�߿�͛]��|]���,W�FAx���_�m 8�����̄wZJw�����l��<�p���v��R�����QR:��8r���ZiC��G�-"xX#T�0�A>e���,�<��!��A��Mm��)}r�e�ś�@Hǲ���c�����J��wxt�7�t"  s�(��>�O����t#a�����aڷ�LA;��ߣ?%]x��U���+($w}X��j]"ق�r�.x (��U3�|���6��l�e}�F�c�0���CmU@�&���C�U6��\8U������s2�ebr>���4�7��mCI�BjX���D��C+>��^��<>� �܊9S(9b�����}u�,�
G���z�X�~�VA�<����l0�|gK��^K,0=���v�~Y<Y���6������/���H��ޤء
T$ߍ�H��*�<R�9$��F��cB�;��ʸX��;2^1�Y���=���`���#���҃�i�p�=꤫�T%�2dyU_����s�L96�
{[P�@US�kx��i��.C����jj�s��f1��2Ib����3�8�?Lf�#GEil�y��=T���f՞-N�y�[Vm�CzFU}3|�K,z��.�v��U4K8@`��z`u?Xga��V{m-Z}þ���\�Ch�+��QI1�������<��D a�f��_�Dנ��ׁ�O����w�'=��i(Yō����1Q�=PvI�ǔ���~s�V���e�5A��Ԧ"����{�2�S���R�x��b ���
�1g��L��x���;jqg�ڸ�	w�E��e�ޭ����̧
"��mA.���Qc�m����U ������ת�U��E�N6MC��3�SH!���g�g�]6ݙ_B4�4Ee��,���c;vn:t�H��Z�V�'�J**���myJ�՗��F��	+�.1m�ʞ����5�0做�$�0���y��1�&��"	�1�#ꐜ{��K!J��@ޅ��û��yV�L����c\,��EG,����}�3���� #r5����8��P�L�c ~����5�/����^���mW�T0q��=���Q��m"�,����NJ�ڟ�#��lp+kQ��Q h�GFL>N\�kD�~�;4A��9�<j�.e�����"y�Bz�Ay��T�P�5��V��� �t��kR]L�c��@L�5Y�MRӷa��w�g�Y�H��E�a��2�H�A�6�R�#�-�`y����u2�ٞ �{G+F�)7 KV�<(�ʵdk�|r7]�x�jt\��s�g�ׁ��y����4Kq�Oy�;J��f�ԇ�n��u�C�2 ��Z;Ќ-mi�������f�]*���~$�({c�~����덫�G6����掵�p���J�"���iL-O;�Y@w������s��9���?4eOU�[v�����t�E�MR�i�w2��&x^S���	~�6f��\�?+.V[���%7N䀧ХT"�b���ű^g�$�_�r�D�+(D-�^҆Θ�H�������u�h�}������ 81������A_���3х^S~P*�h_�n���`̲��}(wYb{�''&�\��茲�|��i�)�"t�=�)�P��F�Ͼw&@t��o���fv��h0{l^�Lȧ?C�Ԇ;q��6�V4�X�3i�x4w�-F�v~Z��0T(�ͦ�s�Åw��_)��z2����&2-c"wǧ���J�Y<F��e�H`�N��X�p!U�dh3��Cv.h������*�n!�U�h������+,f1
N��/��y5�}�5�2k�r��|Ǐ7M0��Phd� G|��,r�_�_�]/q�Fd�[�y��n��^^�@�=~�+xn$'��Օ�+?U�G���C�h��rT� �#��5j�Ns�#�2�1���x����5+!����_������u�&��������|�B�t��������^g@�,��P~���9Ei�o��>�+�6�� ��%�ݗ�0�,�:^�=��
v����9?A�P����T���Ch�~w���Y8@T��<�&��
����@��/"�\f���mm�X��Q��&��Q���r�c�j�Mz���\��ی�<q/G���%�V����X9)!{�����+Wam�_?��p�9~D��qe�R1�0�@کQ`�.��3?b���+uH�-����?Y�*W�<�EMe�ye��K*�����Kv�9VD�Y�ؗ�q��3�������B�r����Ң��\m�+�_]���!�����UPŗ ��{��@s�ң��n��`��*7@����y��[��.��$�Pl��C7T���QN���4Av��ƍi�/9��H���}�e�<��wė�o��?����w��n>�� 3iԧJ�\�����m&�(*�d��R����E.D��Ȥdh�C�E*�yϐ_�2�k��Y��:�(|�*��+qOV���2�w���2�Y`��: #�i�W�If�̏����K O#���?��$w�03o���_Z�o���$�Np	F<�bJ�ѕG�p���ַ+5��-AD��u��A�)��y�!M�M獇jPh����[���-#��o9��Y#��S������&ʯ�jX�bnϥ /#~�Vs��(�=y7#�uX���P��-��]ȼ�(?����n����!�,o��P�!�Fg;Xp�WHIg�zɀ�������� ~����9���N*CK|�ū����pQ�Of��V����0��W�ss�ius�ڕ��R�N#~���U��r�,�U/6��$�k������ ݶ���E�e����f��6�H����4`�VnQ�d�,��%�d#�b��|pl������Gv��/���9���4f5uT�,��<��1ì�]��FS�Bu3��m�ro�S� ���׫��g��g���q�Tw �M(U�k,�L0�%���M^���!"A�b�[�kg�x�l��x��2�ԎE�_|��o��I"R�G�}�5�'��H�9Y�9 ��E���*���B�\b�?��z�����B������L2K�rI�y@���H�Dy�F��+7ؾ���'��$�e�"��A�?���/�����;��m�jk�:b�~����@AU*H,����rk�5a��`W�3 7-/�/a��� �O��̠U]��)����Y�>�����r�9*(
j(�#=����q�@P��G�j]O�4���h��
���W�F��r���(���{��B���B�*k��B�;w�=bl�i'��ާgo�m
W�.���9��������dg$��G���\�?{]8̎�㈤�T��*��y�Y�!w��%�$��B����a��4�������ʔ]��b'�ǵϡ�����tv��d"�����PkƗ���c��Y���:�j�1������Z
7):����D�B�j(���.��wH��H������wq��b&��ޑ@PMS���g�>�g�����6JE@�*r�$ Yݵ�Z�T:4:ۅ��l�en:�;7�p[�F����?�$3��dV4e7��XZ��T�E���";g��� �8%[jJ�1.�}|�𛌽���v�r��I�z�I��	�[��)i�W�Y�]���R�������i���7V`��&E������E+N�t��]�W.$AK�90�^�Ut߂���{k�����'���a��&�������rT�/���hN�b���9�8�L,X/��7$ ��9��)�ƻ�aZn$��)t��Xqo��
i
�o>+�B	I4�5g�H���ryN�B���f\��g��$(d�Z1CU��-P}2�ց4�w -{�(u��_ddk,� �;��M;sV$t��S&(��h����2�	+�A/�N�^�K���H�sN8�u2��}���*�� dz�` �[^~̽�����uCVܘ)&q�f�t�	Y��f�UI���V��b�G�1]�'/�l���&�P�����1֡�W�V7mм0��f�2��'nYMY�,Ғ���.�t8)B�u�:�4�vm���9s��'�NF������]��d��v7�8�fŹQR�R'�b��Wv�E������u��٫������ 7�Z�5�l���rZz�E8�O��rN��/x��؃��%J&�.w�?;����ac.n&5ۋ���:���J���
����X�;��bTX⽽5.~:�T�����/W"��z#�Qyi����ӪK8�-n���05'Ԍ���dC̿xf,��Q�>=-��քϼ�]1O�ߩ��)Wh�d	3�}2�M�����T/���M���>�TK���I~n�q~<�r�^�������s�+OE�N�Ԩ.ޫ�p�j����v�}���d�䘘_] nmyp��Q�w�u�$J�dQ�� �g(>f$+�h#�	`�w��q�O?�T��R1����&Q�}F���_�3����ih�����*�>g�V�o� ���	b<̒��*h&;͍?Q˻���K�m��ܘ�K�@���!� ��	�SL�edb�3��_q���h����ε(!N���P���wq�=���\���8;C�K��Q��W�
G��bgc���M����S4)%��,3�����A1�m��l~!e�첓�ͱ��ւR I-'��	<q�ŐY