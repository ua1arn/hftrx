��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b��%[��$~��0���j����<�S�3�,�%�*�N>��4�5Z14��8���ᶜ~g6�Y8��W
kne�y.-������MʯAF��λ��&��/��eSXa����g��d��& ��x:d[��f�AP/�ѱtk�P��Yq��)���G׷EkkT�s��^����MM��<s{g�$��@a��<J.�����p%��*Dj�wm)ƙ�\s�5�!��"�˿�v-���\n�s8��`��=����\D�c��`|q68OB�Z�ʹʤ�B06l#� �r3����(�Ѝѳ^K�ۣB�P��u�J��a6�V�.B���Lw�.����M|{v|inj͍��~��[��1O��}�>e�h���i���Ss�����Y�\&h��3$��`ҽh���rf:�c�@n:y�dM���\�jT�M{���W���J��Z���Q�	"����4*�T�)>��h"��=�4��5Si�ñ����"�nI�Y7�7Q8�8��"on/9��V�K���6Y�s��Y�*f[�Z���;P����M�O-/�@x��ܜct̠��z��a������`���l<A�d���+ܴ��L����*˗����yS�C�]4���2��1:T]W��M����F����s�c+zVI[`!��(G	�y"��A�d�x9S}GZ}VWM�y�6j��P�O[��p��s��Ǟ[.5�_1�9#%q'*�:�-�4ҞP��a�=���CEU����l�YW�6�_� .�Y<��G���q�+��X��V���Nm� ЗlQz(�Tl�Ai�G�%��s`!e8����]7a��|��>�
�ۚ�@q���=kQ�g�tIt`U��5�jm3d*I��Z[�� �P�v���:���w��͝���BCYɎ6�m���+�7�S١P"�赬��a���O�ᴦ8��-�s�mK���B��#������ٵ�����X_PRd���jۆS��13v��n�V�����h�i�@Ս�8����� �Kj����nu���2bOy��%2��6j�1R\�9�<�MVv�N���#�i����p�A�pd�=�s�y�n��?��j*y��x����Cڗ�uӵ�ps�h����g�柼�����I�u��!3BK�}�^�g�_x嫾�I=O����Cb�F:��P���bQس|�G���w+Kͤ!�?2�S�A�s�<� ;�:uywU�Dm�(&`k�K�4��-d/ݼ -w��#��Ö��],����g���"k�8㆘�����@���Nו���(���:W3���/	�2c�=��	��Mf�=���?��`k�O�-�N.Ų�EBySс �1։G�z���>j��/��X�s �^��R�e4>�h]�>'�s���@����:���HZ|dT�X��+\�`�6��8m�g�>�.����v���~�F�4�׺��)}����Ī<5��/��|TE�u}{�G���9����<�Q���>^����GFf!}���͒�#���h�a��l�Ӽ $�����x��N�6�z�>#e2J���Szwƹ����� ��qa��(��ݣ��rr�OH?Q�ެ��������e�gybT��k"l\���v����V_�;����}�14�ҧ�_Ne]�,���(�����~��1��=b+(P9?�3�H1&��?pG1�K:"��Ys�. N�ns@m��|ʇ��f���i�E���~�	�쁨���$�@5H���8qw�:Ђ�x���'���W,:e��G>�_>�O�~������r=x0j�u���ݨ�(�Рi;#�*�V5.noi����)S3�v���������b�};;�RG��7�-ܙ3�G���T5�L���q��5��daQb�]*یc=9��"���[��w���؝�� �.�+C� e��c �f���5�={�C�$��&�`�0��̑�r��!f�{�ҁ�>��~�Y�j��$��:�\^�͓�02���̋���ηn��ݽ5�vL�*�����S�R����z�+S��8�F\��q9�������_����\T�"�t	3�|ILhHBS��r^��a��n�>bGi=�h�;�6PDI����� e�c��F�tB�r��(�}y��ѥ�F� �|R��99Ov��FOǀ4�K����,,���d�ԉB��i.w�p�?�\��CF�$FH�\�2���8�z4���2_:ff%;��?~�[�"�l�d�J��|~��s���%k��W.�D�s�Mj|-c19}a[~~N�Ĝ���٧�{���j}� ��.���2I�������d� �$���U.{����T�(�a���6��vpb�F�?bAf~��-S!�l�M�����cK4����ߢ�o�4��R����GCɊ(��gt);��gֆ����Aj��J$�U݆(�J��L�>	���N� ����`a��rHOw��o��D���ÊG���P��6��-����G'�|��WR�
�i��	.�P�Y���uV�����1�bV���m���������s\�9K4Q��]�9�9	[��:  f&\�>���[�����N����-8�_U�f�4���.�oT���jA�=��eU��|O@O�����[ ����p0a$a�\�fd��%��y^��}sN�ǘ�[�����ˤ����I�N��}̂��^�R�5��V�*�w�NB�[��:�Z���g<&�7���0� ���~�~���Be�������5���'�I�JG��>��c���'� K8T�m��O'm���'̽�?�-AL��
v�^ʫLP�� ��I��d&t#��T�=�zz������y�
��(����W�#�+��߬����G�h�ô��)8)ET�< g���u�1���fB]f�[ů;��wU8���:�����@�rBB�^����$�%��� �E��Y�4E6���gv�&�x~�2��+r��΍�h<&q���"X|^�j�n�4i��&�L0�]Iɚ)VK�}��J�����m(
��[��3���w���җ����CSŷ %����#��A!���)i����ߤ�����_e:�ҿS1��|��R��TL&b����NQW������֤&�����*&�na�$��G�}����U�:�*�]�i�����C�I$�Ȟ�X���5M�픵���FJ�"g�f����ڊ'Q��9�C�j�QQ�k�̦P�=�k�_�hF�d]�ӹf8O/��%q �Cn�����R�e��vH�F���u�N�g����1�qv�NPH���r�4��3�}�����y��7��u�<K�&�s�q��q�.S�M��_(�~r�t�YUڅ�)x?9��0O�`
DQ�XР!�><�;��JH�������ܾ)=��H4�&#K�
�E�% ��E|��d�J���W�-�|�j�����s�EG���#�U�M��ce�a�fjaD����[�P�F�^%�척��\�Q�x4���o�RK�>>� h�����EV:D��}�Dqj$mZ6/� �4������V�<I�޹��3F�]��8�8@u�v����1L�������9
�.`��W�`궦D#A�q��q{*��*%[/�,��T��[�j3�� $�h�Zy>'�Ƀ$�8]���!�O4r%6�IX>�5���,>V�9�oa��x�:����<��*�/�>�����Hs�H�F� Qgd�)�\�4:R�=���N�4�!����8�EE�U̿�˶;�6񵧰�:�c�e�>/O���f��2�d>c&��� 	��"�x[$B����mtY�Gp�zE6T��^���=d��OC�F$�qj��
������:� R H��f�U�Y�;j'���R�ś���VVҭ�Si���B��Ύ�B��`>��Q�v�)M�l!���E�L-/��T�b��e+�c��R�����b���æB�O�1�bf�����}�P·���4�Xdx���^�FaR ���Mf$��jɝ^���9��Y`6%̅�S���M=E�Ua��g������%1
{͇H{6/L����5U�5�XJ��&G��xv@#�B����O�=����I�l�����2n�� @��j(�`hc�����	"' 8�O�W����o^GY�w��ՙ��WJ��(ng��N�0J:%��վ��睍�s��#<�_�C|D�P�����Ys�%J�P �.� �h&��^�/�sY;)��;��{�g�.i�Pav 3��ۮ	H��T�C��SoGL��	*<�Q�;�ԩ���]#��mۏt'-k�����1M���[�+��Ԧ>�F?{���ֈn�=}��&N@h)MT!hn�eZ�)F�h��F�~tq2{5�\��-l�AWr�������Tf�<�0&�o�a��okq�n�B)=;p�QȵO-P&����.�y�B�Q�\��&���袞J�Qw��������R1J���a<�B���oO�����D�P���`����j���D:g�yj]�E�LHIZ]@� �A��F'R�-B�m�&�M���7�B�7,/��� �;r���APc��$8��9�q�˙99d"~��M�b5G�����'K�����N���&HJ�r�͛��X�%�g�܆A{��U뛰\b^��@�~[�		�Mt�sκ �o���&�g�Fu��t*�6�bŒrc*��Yl���/h����\�Z����*�� �<Mo�8l�i�i�b�Zj�}Xhr�ϧ��:��'=�KY.�����>n�~a�7F;����ğƗ
�󃟱O�_`?�D��˕dQt'Nz�Hq}����h�qC�,�WQ�2��� ���i'��w8=��C��X�*���>B�~�O��DpؚhA���Sl$�[�Pv�Ŏǈ������ߟï��cD��֩Ǉ�0E���I�:BCr������0w��5g�g����~���$��7?2�T�y:��(�H8��MX��3��o��<=�׆6G�B�J��� �/y?��eVnR:E�8�":CC�N�1V����(����wk�.�P�|_%~�r\}�9c�ҚǪ`����-��@ ����p��w�>o�b�N���D����3��O׹l�W6�Se�<̔{��ӟ$8�	���,vjD���g�M���f��Z��+�Gm���k���Er�zN����rB��bjv!��U��Q�4E�S�i��,���m���h��k`1[��	w�X��ת�"�~GF܌4��¨J��v�S��'�� ĹU��/#��ȝ �1IL�z-U���7���#��K�_FXb]z��C�����2�.^!Ǿ��TڸD������(������]X|���c��c��
�g���G��Wߎ�CB������ �n�(��e�X>�+� �]��#���r�Q�,�!y��l:�1kZ�;�B��\��*$��Ku���g8��:��n�]�w3��>�i�̣�v82��I�[��[!�w�S�~� ϰ��.YT��j�h����U����AJ0��0խ|���[���73��4&Qg��B%��!�N(��2+�����T�V�Ҳ'��ѥ�.8@Y��/*dm��ęyT��~�V����2F���U����A���� �L�X���@S�g�x>bԉ�S��5U@���5bw?���r���j��:���4Q��< ��Q̥°:3��L�_>�Z��C�������A	g<���Q�x5������U��R�f�*��>;��B]���]�n;H������H��/�� �Y�ڊT��Y#W�n���z�_���Jy*ϏZ���n�I~U3�+��v��s�>�me�
&��	@e�SI�tzC�p����H��PF�&�s��';9���"Gt��f(���]8P�& �4L�K��1�#�o"Pc�Ah�C��p�CЫ�B��>�ls�G 0E���}\���I��D�'H��N �,ݧ�5��Ckɿ���,$8��e�
(���2�v/[J�fe(�e������\H�����6J=�Z�0���HZ5ph��J�"��v"p��XBz�LKX(�H�:���л
9[?���Yķxh�d���A�������x�ő��'�����!���t���w���R~���˧i����\����	����	��;lXu����dJ�1wܺ��B��H������~��ē-�e:g9���{j��.ND��V����c�jU&�m#n�+F�#Z���L�� ߵ�at$��.�����'�2;*���M��#о��������<�l��B	s�([�0�`�\�B����l\w���:��6of>�_&Kڹ��W,>2�RUN]I��Y�7Ӝ�qӓ4ɂ����[���&��(��k�uZ���d����6ݠ;C�ǭ�!�叧J��A.�,h�0I"u[q7F����������i��*�T3K[�$Xm���D�:�},���\p��-�?�p��vW��ʤE{&"~੬�����X�	='��t�㗟8��mZ� �`tұ�-xc(�&��3N���w����"�\q*X�@�z+�>~[�ţ���Q>
^��-�jzW��1&�<�ysPOIA:��C����@�ͼ��ȹ,�cQݜ���_�ƺ~I%�B˿��R����}�k�!���q���HlL�m�>D��W�>�i0�� ��|��\�THe�=e:�����p�K�R*��Hǔ�p:���-�wR��U�������G����R%,y������&A�`$�0m�n�:���h&�����q�Y7�a'5U.�);P���c>Q�N Pn��ϋ�$y��~Z��DF����?�f1a���Ք1�z�ȱ9[C-��=�mi�d7���B�}Q8���:lҶs�/��Z�����{����S}�x�^]�e������.��;��˟�e@�$�8�ĭW��S��9_Z��8Ľj� n�ٕyΌz�P�5�vrܝ�f���J ���ɚ��y�����Gw"��L���y_v����3�ي����)8& Pn��utd����L�]Ըj+����]�O��K�#Aݻ��[�DV������f�b�r��Q�7�A��D�P!����#>�0�9C�x�7` ��NF]��E����
d'�Y��������H��ۥ3޽=sY��w/��(�+�$]��`ߋV�̩L�M����s���k���	���J�o��)Cf�)1<k���_��Frųo���kOZ1)-��E���dg��-�v$`0�!��K0k����U���/;�"�22�62�4oL?�1�z=
_Β��@�v�sn$�q�o�*$��oti�}\#~A�����N��=ݷ�]�F�̭�.u�>E��U��j�gR#�\�� Jnsy/�-]���~�p$��TF�I�%P��8%ߍ�a�G�]n���A�S�pC��wzv�L`���
�ZD�[�������0y5} JKq��RN�.�c$�W�����iMR���b����	`����|���	{Ye� �YE$X�G+78^�c����?�b7i�`>dF������NP@�s4�캤�&:��@\k��r�Ұ����٧��$ݝ�xj9���U���q�a�g>��w�G~�' �K�l�W���C6ב�쏭����阨�<R\U����\�p
�Q+']Ͻ?_[���u�V�I���H��t��Q��|Gn�������q��Y&@�����T!��p�G�M�E������4y��\�|3�#,K"�c`j3m���	��^�4��\�aO�/��e�S\�A�d���כ[ �2�;ȉ:՞MqU��n*w�(�jA�U$����Q͝Ԣ�q�Y\6�V��=�?��g���ݘ=��j�V�.���%j"���w*C)T �ܒ�j�Q����͐��SL�Ѱ�HX~�)q�=S�a̙I��e)�^���h.Y6θ��fd34��kg�]k��� �{|.���D��2���"ϴśP�WR��
{h�|��[��hK�K�����6gK��h]b�F��|�BvI���p����q+E3zF)���ƞ������nc��U����
(&5;�?(f�H?)���a&Ǩ»iLt[)-a_#m̌<.��1�7L7���@FUf&[\=��b��_��9�s��0T��$���h���(�ugUn�k�\��`ݙ�����d"-�a�jm�Ȑ��Q����~A^���Q�^t8_ᇆ!���ү�湺Dy����p{��8>��E��ʅXK4�%��J��a-� �����t��v��O��}�]%��P�cM��T��gu�sDbJS��k(#������$
���bB��U���t,�,L0bT,RK ���dͯϜ4q��n��Vv�����]�͢�8�}�$������;���'BxOP�^ީI�8j����FEr*����G��&�'��͓�*1���������;a��wk���fq������|��`��j�*O�94$V���?��/I$�&ƻ��s�(5��U9J�oɭ%p���Ntn�����:�D����nU)�U�U-̆�ɢt�сn%��bn�e�i�����ɻ�2�"�Ŷ����Sv��o�׼�(q{0E�����{*������~隹H�Hzh���@��M��
H� �vi�ё��Դ�LH��[�-�^B�Ixnل��t�����	G�-�aUE�����|���`f��=Y>"�)6����ë�Ȟ}c�������������A�e�5W:��]��$���3&�-"2P���Z�P �-��\A��t�Z-��Q ��%���:n �����/k�+�����kd�ޝ�PX����W[��X)v-d��Ж�ZL*�m6_ ݰ�Ԇ:z(e�6IV�Q>�~w��j�"ቺD[,�C��꫊���(p} l3P�SrL2�8��§�ؾ��MwC��y]���%���:�ѯ#��C���j.��ۯ���xٻ��ŲW�ܵ�aj���L������µ$�0b�����6,-P�<�,���;�P��t��7�3�����N�c��C��.7>�}�WZD@��;��2���񞞪?���n���@
^�:��<k�_�>�eMף�U�O�V�E*>������s7*���'�cx�8��ݤ���B%��7*�	Y��\�皐�3�iK�mid6x�H�*{��J��y;�����������M���R���?}-�Ua�<J��� �BY��~Ӵ��R��AM��eJ�r<jF�JJҐv��P�E�	��3�^uu���ߕ�Pr*;)��VJ�3���M.dav���R�y-��P� �L����Zu`AqH eU�\�vsh�j��0�GId<[�����r�P`�'�h�'�M�� ����2��b/��j����������~����[����
���/K��xf�6q������c����?�����X8#ͽb��[;�>�cϘ� ��T��&}�8����a+�,С��7ԩ�5�J����
�&���`s>��6'}�Zu����~]l�^������*a��<���b���J-qP��7*Ҫ�Vq�# 7J�D[�:nii�n�y졻��r�����r�c��Z۪L�Y��"Ƥ���������.�j�����T��e�]�y�E����&QU�&��t�Z	@���֍��dm7zL���e��)�XF��$���n��	��1���L�y2Jww��I�U5�uf"��^R�S����\wu��7TΪ�=�e�I�ۧ�8==ѯ�N�^�)F����Ec�Z%���Zi�0`������{*?��+Y����'ކ��w1�N��<�e�k��34�1�6�۵%Qh������=���}�;ռ7�rA���2G2�]L^f�R{R�����C�:Z���׀�I2��0Y����Z3M�{��s���	�A���JԀ�j�w��ͺ�\mT�1[��E1M=�*��~f_�˂	��k�����2K`ݜ2��p-^��O�`1dJ�8�J�Jᮮ��崨䱰���5'<`��n aRU3e�t���������P陭�q�����dք}���k�$+�ҭȀ���u>��%N�@c�`>��S�CEI���
7�������[uXq�!�ޞO��p�)�.$iY���	$���>����z���y���"�DOqө�U��ˏR�eRz�T��(��o�}n<2�M K��{�w��u`pߐ��6(bpS�\u�8&\xP|~�8�
v�U}�A�cS���l��0��x�*(�R�jQ�_�"����4@���3S��]ԁ��=O�a�/�F����L����?�n�uc&*���¯ݷN��^�@�8g{~��JF#����R�^N��ކe_Z2O���w͉�t*�m�H�x�.,'@t�GQ�ke#%ȳ^�!|��Y�K�"���4��,����9w�^��`���Sc��Cn����qG6��9���A4Wփq�+�|ն7�8H�%&|Ps3�GN2L>�*�tr��(B�n�M&���2Ỉ^��\Ywϔ���4w��`��P$~����I�3zV��QVȵ'��G�Ia7��Z�H�ҫ��{�(�����֭fd`%�e%�aW��#���x\ @p���������o�5'����Ѓua�P��`��S��)U��NA|ȢK���yPK���!q�:G.!��H���Vޣ:#�Jo�S��|}� ��� BQM�*�Rf�
ZxNY������~ƙ��-�M�АG��"���}@�=$��X 	es�q��-�_Zl�´�A1o_j�#�l������h]�`�ϢXA:l�ي��ڛ�9���e�FX�8�N�[�>��OdE�]��؁��CPs���?_I�/���9��e��chR;��P��2+�*i�>���u�>���n�jz��p��X3eԟ�k�E��s,3d���t|�4+x��q�ͽ�L���Y���:��w�X��ѯ��HD%.d�w{���%֥�oa�x�HWp"��J��-8a���N��M���3v�U�Ä]ͪKO쉂��Fbl*�ZW&�*�$,x�˒0��b�i'�2�a�SO3�(L� ��<c�8KSA��~L��5{%*G���H�Y��MKm�r��n�8��;��w�u��8�I��
�7/.��6,/n���� `P6)�{m)����Jr����_Ȭ�xM�s��1튊�{���}�&`�<G.�z�`�c�;��̀­��-�����3���?���y�1%�x&dQѢ��>��郼��ꓠ��'G��v�O��O&� ��h���Q�"%u��!����/Ǐg������x�<���y�!m��G�u� ���uڒN6h���u�	]w�B�Q:��+Z�1J�I ���yd���7a��i���a�9��¿*u�?iqzd��=c�K�̣�b�e���	u~���A��a�`nZGkJ��S��� �q�#C��2�1Nz��}V[?���~Q�f�ܺ8�4���㺃i�C
{�үe���cӟs�C�ʭs!�|���Eh����q�["�	W3$3<���%�^r�}k���c5u
��ǮW�����Bj�u�E'��bUzBA���n� �,�T�j�r5s?ԟ�Tr����"�t4�p��,˯�=���������#��1c�e1�`���g׬=�����V�fdL�8�|B�"@��-�Š������8f�����yd���2��v���-��8��Kx�����ĝ�|~u�
J��3�	9��l��8�hZ6�CY�d��� ���i�8.��l� (�z�	k XHc5��HX0�����,��>�ux)qh��̊C;ZiX`�`��� $m��l�>#���%C�'���a}���꟥wEk=�>sO�&��0rJ��s� �ŀz��o3�<KdyP_�����P��9 ��*��1�MZ�,�hv<���Edũ3�F��,C?�	T�C������E޻Kb�z<��_?t
�C�Y� �O����蟮�Hr�	@D��N�"f��*�ᰣ�2+[�y=�]�<�G���I�AY+`9q�w��n�9 �Jw
�6r�E�`�j������H.�� ��=<"��ó��N)��K��τ"��ޚ�9�&�	��.bgS�,�i������A�ڄN�C�nf�7�Н3)\�0m�F�s+���4a�~j������D��ZCXK�{�=���~K�W�l4�p��mFf�)�}�� �pв�:��.��V�[���f��!�_sc�x�y:�%�&�g�B��9{¢�_r$M�2EHy.�u~�y��s��A6���2��0,I��W67v�< C�)�&k�!�8�Ѡd%(!(Bɇ�y]oSX=%��R�%˽>�n�y�ŷHG��d W�玄z�3:��]�Id������-�!����Q#�~0Il�̧q���GV@f��J>�|�Tc�� ��h=)�D����S�򔪞Z����8C�wW<[-�&��t�'F߭���屃vv����>�+\<�pG���Ժ�U#�� ��rȷR��f��t9.��s������c",dm�!'��~��0��AH��O�����.��4w�4G��OG\?�݉5���?�Ⱥ������E�C!��X�LW�*���E��ۆ�B�����5�R�x����pʦ�kQZ�k��MP�寽$����1ҽm͠/�R��HЬL��Etu'«�p̈́P���=HPK�C?�Gb��,_ELo�0�@��cL��3�bi���|f�o�r��	����ҏ�)l���BPz!�@²�S~�Kx2*9h������fTTe�`+���4@����1B̰��u*�����8oEby�I���q47�k�6�a�2H�@l��=ϕ�c����u�>�
������c����gfj��Ϡo~[�K�K�$p�P��E(�-��^2���j��,׭�v�R$H�р��O�F�B�u'%ف�Z�����I�|�~Ǎ�.�4�V�-:���O��]+���y�Ƌ살�-	0D�^zZ����ۄ�U=f!�Αб�Q.�MȼT�T'b�� ���i�ǔ֛ps��f<{��V�t��L�g�6#�D���9����H�r�a�g��q���~Gq��߃c}��7
Zy�\��z��� 4��ӆ��t�\1P���j��gܵ��Lɞ�-5��1���-�EUdBD{�Z�]9a#�4�/�tЛ�=O3f��/HVZ�����@8�)�76��l55�~�A�A����}�w�?+ ��կy.���PcC5��c�U�7��x��t<�cUÒ\߃3o�w��셳5��Q��C5�R��{\.���H��8h��9@�?Z�o�<��x�r�Tg�t�w⛮H#�o��u�"�Ԃ	��
 rOk�ơ��gNx[�յ�PD� �;*^N5��~�@mH�e2?��ݭ�Xy<P�V(�$��\�+c�K�0\}�,`{V4C�f�5"[e��^��5���c��v\8���}p
H��P�B֭q�d�|y��=@�w�aKB0�M�l�/��cR|f�����7b6�>}��Z! n�,%j���m��+YL�NC?=�駈u�8����$l]>1�j� )�+X�9Y�2y�i���Q�QA׾��ff��j��D7}�8e��?rF��0 �)���'����e��h"�����zG�T԰���C�b���N�j���-�'�3E��vbҔ�����y�̼$���b����Xs����o�[�iD��U����R�����G6��zVO�%D<�Fg��-uԼ���k��d���#1Fc�{Fo)�o�X^�%C�r�E;@�� %F)���L��1_� ��� j&|��ĭ�ur'19�&�`�JM� K�,BtA���ى����ڸDu2�BM<h�`�A�lA�<tu�ͻ����<+�@� ��)��es��������.T��Ћ�u��X ϴ�H����*�����,�\B+��0���:��!\RϽy�-�E�`�p�~���H ����BL�w	HUw�$����������΄��;���Z��������8�~�p����[<Nw��t=�m���&3���(��=*����4���MfO9z�|���y(*A#=\_���ؿ,'.��a�HY����>�5.��<��&��-5W�΁XL�{g6�혴C���&�,�m�n��-�����W:���܉��<,�����J���(;��ZR��*o�|rk�X1�:�t�:�x'$I�}Dh�VJY���[(x:t��;}�;K�S��m*��r�K��--�B�,��M��-(�N���>`,=��Bl�\�	s�����ǞcF�2�'/�(	A6Fp�<����Dޅ���O�w@*�U1y5�Skn�y��e��Gח����a�:�S� S�ڝ�9��?/��x2D}]9�~��{��/mj0�Q)6]G������S��SW�ڠ���b�ZH��&�����X˓�U�)X��)x9�����5૜(��5�Ğ�7R���V���/���t3kF�Az�uQG��������;Gr[�*tB)���n��.�fΞqC��	�H�^^RZ�'��d�-]Ң�>@���U��n(qġ��y�S�e��pf��0�6]����-��"�,i�?�І����Ǔ]k�Ԑ�%��i\�)�ye���R؁��fM��I�q��(5�i�eLF��ek @D��B��u�_)�NM���
��G�?���eU���\=�}?������E;3�
�^?�[aR����Y��W��N�R�sB��Zq\p� X�?)��Au��a�[ȏ�>
K�t�@R���G��K��o�� ._ItT��kp"]M;�����"󩣆�mi�>���~��'l��fՉO�L'D?7��5:jP.�='V���;�[\Z�˩��ِ'�֚��VKU��]�!37�͊�x��"����(sپV�<:�F3�U�%pEw�Q�_�n��U�_w��� �ؓ�b⨰R���9G�m^�S�,T�ZZ�O��7�yq��4v��9,�aYȋl
���U�Z���q���)j�[Q-W5Ã��8Oe�49o�*&6�Y栐����9�ʫg�Y|ٷbe��QAf���ܵ�Y ��&���v�>�7�$�*�LQ�y��a� �%�I�%Vp-m��BӃ�a���t�X��|r!)�}iϸ��?�
�ȅ>���˛�����e�@k�b�EF?[Dj��W�CS{2��E�TK�T/�װ�o:�a� ��7�^��2��s���~�L���w)����T��5<�~��B���I xիX3��-�rv�q��m���o��2Kj:�G�Mr�tI����~��s0y�N2[Y �H������p��>ER���RRA��������A�u<�7rlI{J�
�!1�,��	{�.���D�`���eA��6F!����)ܢG���3�d�7�-
PRJ���4p#��G޳�[-��"\��{	�$����<X ի1�R&���p�
=��7z�G�g��:7����U��9�+�bB}�G�S�V,':3wu;u�<��V�q���(a������z�(���ʞ϶���3���윺[T��)ua�H�"�����ϭ��2�'"suт4-�͚A���{B�a
l}�iG$�^,C�yH��N��1P�W)�7����� i�T��-.�Z��?����7�$l��_\'�}<zB�p]#��kH�M��;�ҹ��O�8�lI*�	���a5�����nq dYtəb��A��
X�T_�����y;Q�)� �q`=��ER#Wt�&�B/��u�i�q#�/\�B����(2��d�p P�?�]P���Ⱦ��d�L�����QQ�ؼbM��LA�2d�-��)��MXO`@u]��<˅�qn|�&�Uf�`V��S�mOȕ�f'kA�ʼїŞ�j Gx�8�m�ss�`�;'��\�r�y��%���5WoG׫��_��Sn�-B�e�W3ޤ�#�$�OL�R��3�}�ap!c����MQfNi�|��n�U��3O �T81�9<M�e������?�m��}Uv�d�9�h���������5i�YWA`�Q�1���Dl�H�Pt"�Ow����ߺw��i&�G�1i�"�(}�3��:h�O��Z�aQ��7����d^C�i�_�?���}���	��1P�ݲ����_���K���Ϡe�</�i����P�������{�>�蘳���D%{	��I#G�|�����{�O�q��@�guBs����f`
�!�Ðz��&0���������to��"�!�DZ> ���'��徿������Lٌ?�a��<s��c���I�j��pcX\P�h�O5٢Pd*#丞pҦ������'v� h��*�N�������z�r��l� �ڛ-��M�0�~��KcPt�e��-NB�2mE��"�"_�
v�x-��%Y�sne�n��21 ��I���#��Μ 3�=\<?~���nB��_�>����#���̓�J��%�Ρ�x����T��l%r'>��uer�_������oj�ƍ�Eg�������HL&'���W�Hc�>�b�"��c�⺿`;1���y�5���N�"�1��z�W�p�w��+V�u=�GA4��������OU��3��m�A���#��@�8U��D��i�߉u����/>�O-Kd�h |���)U֘q�|)4H���TS��XPh��Tjf��;/���ہb�?�����(�L>�6-)�{��	�[�I3����hJ�((��$��G�j�o'{t�v�7���7s ��9�^.�����	��6آ �O
ڤ?�)%0�-��s��o�����-{l@�2�����*�׵�-kfaػX��%���8�B�b~y�|Xa�U �R�{x�����z��~�,<�|7�I��w.����Cs����Q�E���{!$�P���Ch��GHG�u��F�|�V��ӭB�>4j?�I×���G�Hg_�@���'�3��'�����(����Syeˤ��O�4��,��c�"� �&����p4�,'|�֝^F4f$��L�v5>A!A�.��	]l�a���H����P/�7X����G-�u�B?��"�f�XS��B��|Q;Jܡ�K�����.��^Q�Z�˗l;��a���A\B���M�d^��dC�����B�ʦ�%�n�+-1_�Q�hf�0g�����\��e>��fp��sX�n��$Zi{�6��	�K�^�X�j-^���"t�gg�i��4A�T5�pK���z(c�����ݠ�m���J�����<����.�6�Cn�Q?�ǨۇxF�x���6�Ou��sHb�
0�|R9�< fe�����fe�XSa%
Zކ"2���z@b����+a�?wQ'�e?ܵ1�*I!l<�ļ@2H!5e��j���-hKą�L��&����5��z=X�i�K�W����EI��p�u���7�;���O�M�;�O5T�����]cIO��A�A#�<4���#�������<�2֭�E3�!��"����]o�T�z9�D�saE�yFeז�oj?C�`�(%&,���M�%�Gws�-����S\��+�1�Ȓ:+���[X(��\��g�v/���b��:��g��Z��㸦�+�}����CΘ�^Zsj�,�N��I�?������,0�*>��}�ܙ3���L���OPs�m,~d݁�Hcz�rӑ���]<�~�� ��Q����*��/9d���:"�ߝH��l�� ��\K��]���L���0i�����ּp��9���9Xt�ݶr�Y_�� &�H.{��wV��Nd���ƾ�WF����/�W��w2 J/�Q��YxҐ�G�������r���OU՝��k$�$EMn٣{(Eaw*_o7�kN�`m*�Ó��$�Z��.)�퇅�kPH90�O*׎E��M�$U��9S��7����D'�f
X 6y��n��
�]�{�II����VD��m�\�c���^��kk��P(Q=��&IY!��eǌ�>�ё*�L8����a!���C�Xڝ R#�_#wuS����<z��T(Y�X�DrJ��N�%�Z�V���;�n7@�u�D��,$bѵ�}˽=X�y���eH��;�'���nm����(�(����&ax��v��q�]�G�`>dUғ�x�S'���2�������J��=�b�j�%?�)��=a[�h�Y��_� �p�'���(���p�zZ��Ϣ�]�$Z�M*w�a�]��_8=Q��a�G�>H��$�:�J��J@��A3]��MR�UL�ʗMSb6��y�|�Mv�-1G\�C�.� �>�g5�+���q>��X��*�{4�{"ڿ�W�v����U�	�FY� 5E�i���@o�<ҶV��
��I�Q��w�Ϯ�?ݬ���4/�����S�E�	�?sY��"����J��ĕό���¼;>���L��~��(f���W[۰�NS����n�e�����rA��1��"VuJxǫ�>��uG���gʨ����x���jJ��#	��SB�g(_���f��R���k!4lyT�-��`�#���tH���{>=���F[9����Qd�>h��a�^7�E�
Tq��wN��;:���8v�4�e^)��ڳe�9�Y}���@���v3�wYب;�� �E�v�
�w������|*� �X�އ��ӵ��5��:��c�$m�c�ch�ڐ'!r"�w�XzP�Qg��7�W�����)ߛUT�y����!�tU��h��d/7V�8�����C׏Sk��vܔ�.K,:�p�Y`�*��4��+��c�e��p!Q��g��k�	PNݫ�B��5�����.�k X������g9��|{�m��;9���#F]b]�]h]2ȆEl���jSf�d�v����03�p���&�DO�\���!qI��娹��Rph�(Yid2�����������XT:��@�'�a��]�o��ݳ���zgx��.��Y	h�����Sx���e�/s���+Ӊ=ž{|w^��yE�V��F��C;����}ݖ�r�ya��� vh>�`=��-P\]b�`e���3g`?�6�ǔ�'��p���n�3�|�jb���!����ؖ�J�w�3O����砯�r�o&
"��l�F�����m�r�Z���=�s���R�;��k�6M�r��t5����y���yY�[���ؾ�?�Opp����������.#�:;IS�S���#��|G{ݽKS��5��Yn�[�4Z.C�d�\�7��qj�R)��P[�5��߱�T���=k��GYO�@�/
�E0��h�����-«#	�yߨG�T��
�I1�iH�o��O6
 `SGgOv���š$<�Σz�AQ!M�K�~�1V�xAF��"��ʦr:��b��kʖ*������6���]Nl����
M�|���J1\��*�Zm�&��H��7E��ܥ����x�壖���Ng�<���[�#����d/e_�yA�w��o��:L����h>î�"�� EΒ��O�
p��I�R�C����W>K����p,�ܠG#��'�^�s:t����-o���j�����,�1�e5ʱq����>�It�4g�N0)�{�
�$��"W�7�;B��'��{ϣ<�F\�rZ����U�J�\4������U�2��/�B�Z3��g�@����&Q0��YJ�s_�w{I���Y>���EA���������"�6KR��
V6sw����*;���|5�JzT�z�i����,����Agmؒ�۪:�����k��[o�O�:T����*�`�u��ƄV����w?�",�lZ����8y=6�tt��O��A<��t���f~�%��\ܗ�lx�:�/��Jb�Kv������ "#���э��U Kx�򷡣��1j(��nBo�fl�s3��a|e�MV�(�j2��b�ڟu���:��ZMw�2W��/���š�`��a�Hv%��m�����ҟ)�5��� ��'کY}؝��S���a�u���3��:�w`D��p7�3HO�{�vQ�d�׌���R�2W�[rH�* g��jk�8v^AA|y�U�������-�*��mE���+bC�|`>����c�i�����"���gn�xǰ}�*�i��]���XFGdi@$����P�y������+��2�H�MkN;�Y�4���C�*���[*G0���[;�0�ΩjQj�}�{��/=���S�ج&(��jt�(εʳ�[��9|I���O�U�� �SG}z퀁�("��6�Z6�=��-����Z�GV�|�B��V`~��� ��&g���s:�uv�	H;V��.�����~�H�|S�'�	��j�>�&�S���e�F���'{�<�/K0�g� �}��xPɷ�H�W8�x�ԚC����
^�����;m�s�4��>�
fh4��	~����]�~��l�����Q�c�{�2�}��Q�}}�nI�H��#�g�y~'��[s����Tێ��tUB��&1�)M��.2$�F��w�ueɄ_�%��Z���x]۸��?��x�:W�܃���
����}�fk���N� ��L���j-=(��JD��D�s��.LamP�dH1e5ފ��^�-M% Vu�"��H D�������;>� G^J�？-�{E��E''d�:�C�ŏ!�MB���I��aDV�i����{���;�����Q�Q��Y��"���یt���*�j�<�>��t��=��5�ɓ���\{Ć�w��7��n��г>��%s���W+m���W��_�2lf�b�U��K��$��&�<�Oz?�"8�|T��7Y��*FV���إ������J��=�����J�e�V�N%�|L�'�����:�E"��&���(^NXxR��i��������/rf�ކu�a�K�.ͱ��mh���/��c3����O!�Y�/1D���G�*
����`��ᄮP�g����/�k�+�f���]��Q�Y��X�ֽ9�;8�	�4�}��l�
�Ɔ��U�mӺk��yKH"�i�i��7CS��G��S�권�A%����e����YgX��q2��u��`�|�|��?�ˮz6��ǵ��a�����`�W��S���
��+���/��U�⒜fx�z�u�|��#�e�|J�w�*i�`K3D�9�?	�L���/R�n�������CK�4���̍ ���~��C6:�J0Ό�;��#~�|Mk׷�J�>Υ>"@sO^�"�7�&���jQTn]�~|:����	�#����%�m��C���G�eZmYs˂*y�I���9��8~%��K�ev����v۝��]J��R�����RR�ɥh���ÿ%�����Q1�~X(�c;�A��:��JV�]Y9K%�����I=ҡ�Y�+aəEר�iTw���O]���M$�w��j1}����������U���&��{dDf&x�
Ʉ���a:����]_�qV�͚�D����&
q�c����ʡ��Ҷu������5�~�6�:*�(��fs3�J�H.Ѧ�P���F�J�l�ְN���x
�44�u���1nh�ǣ�TY#X<�a����A���_vo�kŲx�D����V,j��dVvh)��ײf�ܼ��)�����{�%�Ӵ_�Vo.��a�I
���L
�?����#�6G\�ȃ�{�����dͭ{�)����Ei��]*S�H�9M�*A0E���ϳ��|/�]��d"��g�a�,^A]a��Gڔ�f��
oa����ѥ?G�7��e7�R[QF�f�2�o����s*������0`��~���B��� �8�\�,9�jA�Q�kA�!F���_�钻T�&�j���kE"Q�Ms``7 �
TY��|BC��ͯqQ���-٫El����QB�H��Y�ON�BO�����c$ڂE�iq륈���{r��*�	z1U���(gsW�T�>�ǲ���	�M?�f�5rDҤ�\��X�HC�Tdal�����*���r�c3�h�p��Rd�Fΐ�5����*��2d���߫�W-hE �V��Ȳ/#p�+��'�3���4�5& �|H��e<+��e��dON^������G��
J�D>�P�WOu0�:=�/ji�jLM�?ޗAt�p���&�/�1�ӣ0=��y\�Sc�;���?��D�|��K�h��C��FP�4�����k�(�^�F	:_<�FU�`��������r�lcI�c����F|0��E� �Ol�% d+
�n����4+ 
Ȗ���hJ0����Y����бl*���ޢ�� �^3���|����@7��X�Ô>�4DIճ,��J��B�ɦ�7��7;
Jǂn�q60��|2��}��%cޙ@i[�<w�`�t�����b���/a
)m��y@tR���`z:'o-K�D�O����%�q�z�p�(o7�*kY��(�J����O�"��sHN`�?�'����e�>�����1a���������3����51�F�!W�p/h4�ß}�.��-��ZFf$���S܈�)cW�x%S�ܮ�Z<��(�Ê�f��$'�L�8�H�!E^��]%ma�����Fpsz�O��(+̣�K�gq0vm�xK�|�N�b��l\K�'���%��hdY�״��m��gK8T���vF`�l��a}��؊,��R�=�K�	kă]���/��MMw�G��Ά_�{bXI:Nup�S�-����q��/������z�d����C[4;Ki
 t���3MZ�C@_|�b:�+�&�Z���W����(]��trf������^ }��m�' ��ַ{fƪ'0 �	B��:��~��w��r����ʳ4do<�<N�O���*������X@kR l�n���H�	6sx��]#X�Lq٠�(浰 ?�&��*\��.-�oHΦ�ქ��0��˺<ht��g��FS�_F��b�o��|�X�Qu�R P^� Mlێfm��h0�:�"A噬�*y �nwla��o�U=i�6����6���{�bh5�qd4y��8�r�>�N����jt�����G��B3�q`<>+.Xe��0��	⹱�k�9f�M�ÿͻ��z�k$�ӵ�k��MU��O��.�Zc&E.��$j��:ؖ�a�uT�t��k ����~~�ֹ(J1
�|���\���j)r�ⵧd�j�˼�AB����}���s	�vg|�
¹���7u�#���/�k�J��y����8�b�*o ˣi#[�%�5�(����\=����g��V�QX�|J!G�:�Xd�%�4k�LD����]�_:���eAw��%� V,��ԣ�E�1���$�V���1���J�u�+p��GE�mW|�eʶɞ�c��[ 5��R�~�ɐl�Ǡ���,Wi��Z=켻���gb��[�1��bɱd���װ[�!G�F3#�Nh��u���x�<ho��m4*�Zh(3��J�c�u&p*cR. l�����5q,k����W6Ґ�w�V#�:'���l��=��_1�.౏����T��u@2,h��4�����i�����T� ��E��l����u}�}+�H��Tg0��iFku�*����@\����#����-#�Ǖ��e�R�Of��e�0���\c�A�ɞ�q[
�w�S���k�!=g�&ec���$�V�'�z�ma'0^eo���Of����L����^��1<;C��,MH.�Y��Oe7�1k�X�5E�c�b-��{�ŕ>kV���
Ϋh~�~OV�h�)\����>��+TT)���w�=%�G�T1�L���r3�d֮�|��p.�*c�!�oS��Ä���ݟV�Q�	���t�e�?/wfk��4��ˉź�IeoE5Y7;��<�U����XC�s���T�.�.�GR&;�{>�n��?��@��W��x��ɶ�,��ʔH��QJW�<�{Ĭ�ЎђG}�B�q���F�Q�~���fG����|�ݐ?���_X�`��$�V���K�T��g��|Hh`������e��m8*�6ć����o���AHs$���.̙#<X'�[�<m�w'|�{��}�����M@Z����֍�ʷ��_�\�J�ާ(v����8����ZEF;�bt�r��]T� ,��''\8h��G����t7�:�
�&��%�ǾX�kWF�G���~�my
�AѳӇ���Q�w/�KkP��>]�����q/_OU��g"��>$$� �B����[��?u'���㰲������*E��������,H95+TRƥ�!i��c9R�j��h
��̿�J�^�g����>Up�r
�1�x���+���Ǣ7�GV!���E��H�,:n,~��>�� -� �Q�j�e��g<�a�����W�_�~3�d�ĩL�[]�b���Xӡ�%>����)��l^�]Qb���_?y}i�4�I/�զb��iO�Kx*&YҤ�1�*�(�yi�Ke/a�0b�I'�Q�
��-�"�'�v?{:�/˶�o��~�ԗ:���k봔��_��I��$�tN�v�S�}^	�tyx�$�'��Y&���Sj�_ڲ~@�̴~տ���䥬����N�Z�ˮsΦ�B�S`��Υ~�A!$.��o����`�O���y��ʿ�G��^&d+���B����z�E�D�P~,�p.�1)�=G��1�2D�(B{�ؚW�p1��/m�����*���_Z>������Q�	��C��0&�qP�N�ׯB��>s;�T��I�;���р~T�ށ��7hPk]�!�)�I�ZP����hu�fg�4��!��ؠ	����sM�%�i�(�L[�Ԡǫ�>�!C�S��F�w���)%�*'����H���]���,m8�����y"՜4k��������t�MҔ�A0���x{���*��vdf.\v�����C7�C4��k�����*�@�-�� #mȘKwM�r5��]�M��3B������_����_ZڒԜZ���-m�:�L�]���zh�E
��>�Sj���ma�
���ы�R�($Nc�U�ڏ�K�����A��Ӆ�W�����?�յ�y�y���A������Y9^���gc��$qv�GIn�����/>���G�y3Y�'�>�Y�Ȓ\�E�9L����	\�V��o8��q1+yf�ţ��b���O�&��Ɇq�֞��/�kT���Uh�i�z��S�y���K2�ȕ��r?��a˻4PrB\UO؜UQ�