��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+��mHflx�P�-���|S$��R�#p����b^^�]��6�~�M~v\'E{���i M=��&�J� 2�<�0����m٘�;���Q:�����z�w��QT��*�d�F�����05��Q�Kz���g�k*=�M��m�%+1/6��;)O/*��3���������0�
2�V�����Zx��QӮ����E�J�EpEm��^� �V�.8��Y`kT�U���B$)�h9f���<�7%9�P��Q�ۊW�p��i����o�
A�h��MQ�&1n���,�j�Zp$�(�	d�N�]
��f�Բ�=�gCo(�����8�I����N]Š�+V�}��=���Hi�~t��!V� �~������^=[KL�<��* �F�W[��>0>��K>��o����":5=�����&�V�4Mn	��Rn���c��I��軕����9c�[4�4A|n�E�����tRah�	��>���sĄ�+p�n~��[�@]D�'*��:�A2gōt��-G�P���s��q��wl��C����[�������pg��?���r�=���a&B ���V�j���7�r.�u�l[Q�`0�JC=I��%bC.r_��'�mghq.�v� ��nE��,�~?ʫ�mI5��%�5P��c�@	�)KQz/k`��Ǿ�R "UTc��JmwH+e	��I��Ac�y�[�>��V~w�`�鏝冑1/�����E���t��ф~63�R��#�qݳ{�ħ�&����oJt	�����$qCԋ����Z���!������C�}o�7�����V�t�~�Ș�U��]P��ړ��V
���vP��8��R����=ypX	�i�o�x�r����[MCV�oQ�q]�농���V���P>��v�^���9D=I�ynvP$]���_�]ګisO��2�Օ	q��������e?�\6���	��r)����>�*���y`۞2�����h����.�Jh,6s�l;�����}��rB?)���E/��'cZ����H;�Y�~�|�Q�\�'+�-�.�Dj@��%��f逋Y����zs�Ԝ��?��$�3#w���K�&zM�L�G�EU5&�
A�ט�מ���hme@#���#ݝV���X��Y�(�g[�HL5|���Zm�2�U�t��م��2҆�Q�sN8Y�������T
H�Co�`�����eL����Px��A�,���
�<�Ev~GW��0n�M4�0���3�T�*��{�W�*�h]g6���^�^��F��M̘�B#!�1L�Z�&Z�)���p!u�m��$�-R�HL�-<�j����HFM �(mC�s����� ��!���ku,E���P�vv���1�I�e�#U����iJ�d�ʋ�aXb�����L����TX'|\�x������U�u/�q(�G*� ��:�����AM�#��&#��@$$�T4���c�&$~�8ʩ*T�m�c�`��񐳜� �u�b
�Q\i�N�F��R(cia ��3�E�£)4�Â�.���g��i	��[*ѳL�V�Nb��Kb�Ϡ3�v>C�i!v ��3�-�&��\k�Bn`�?�������°]��&(`V�K�´<�O��B?�I�*�g���1%źʎ����#dX�fWJ���M$�X���܏��2+_�˒Qg:�mX#S92�.`��es��z�	�>�Q��ᩒ����&��KzFD��?� ��Pg���V�rN�'ҽ���D��6q�щ2���$9�(�nɔ_����y<�;ba�ß�!���,G�D֪�Y��$j����4m�\���.կ0*%x^�o>?7��J+Æ=����
�g��I�c�plg���|1$(�	Z; '\�[���(��I���ZG�}�?�2W�2�l
�-qtG��d1 L̚��dU�*�͜�������!%LY]��Ԉ�Z��J��q$hNɅ,����� �^kU{w�*e\'1�#"�'��.KԧPL3$W�u´���)ٸI?��EsYn�P�g1��agܽ��Q���}&�����KH�K�ع���҃�����h�ț��&��]B�xb�≤W��K�|�=�J߄�]���/�?2z�	|ZC�Qβ(�!��^��䳂������2��	&N��
"v���f#t�j��BO��(�a�ˏ�&,�%�R����v,e�kfZ.�일�V^���d���E#X�e��M��O\o��C	7�Jf�{��(�}�B>���m0��a}te�CU����(�R��������'v:�;ؓ��h�Ai\��l0]+-W-�k�xD}:q�g�Ն�@��S�Ӌ�Yx�q<y@i���-Gy2Fr���)�h��3�x3u�o��y^� �o�T���V�gҡ�	SSn�q���PV�	ѥ�#īw�"�<��2�^�r�W������$�DNv���e�����oN�� ��F���ί��σ�t�L,��e�&�p�E-L��h7T[��T�޹�22RtM&��#��ie�C�T�Q����E�Q�K�q�4/�VUg7�kG���k��I�z�V��x��2 w8�,\��Z8!?����w�eӕ��N����F��#(j'���6mv��{'��0XK��W)h#����tAn��G%�`�٦��!x�V�F.]|gC>g���<S$�}�[�<�a�<������*�����<Q)O���2���*ڽ�k#{q�4 �O�	Ex4کOz�Va�)e�l]˞�鍡s
X0�9&n$��mJ3�}�����O�Z%,-,��4�_<	�c�V
&�O6ݞ�M%�(r�6���K�vn�!�!�y&�^o��[S��!�G�����60�A�L��Ȑ�ˑ����s�x ������E�j�֜G�S�׆�@w!P�hJ���� ��,nt0����|cP�|��!R{���ޟ4��B��,=:`<��,?�lW�7sA�����o�u����.�v=�{����_�'8�����$��u�4T����vȖ��ǧ�<���G�S�Kٝ
d��}	䉥xVYN�c7��ط������_�v^^��˙�~N{�!�=���3���S�oU:g���%�n�)y���Я�+��Ǟ�/|;�_���s��X !J�]�p�'k����0�o,^1P�g=����u �ߟh��m�8נ�K�=�+�q����ז0��z�`S��R�e��g]0
k�Qb��9��2���G+ks���5�Zw6��._�%γƟiQ!��I�EI,��S�&�Z�n����6(ٸ�T�X�s�r�|~�B��!����n��P���C�=[Z&k�e �(%;Pc����YB�ٕ����o�V�|Z�+-b�*�aT���Ğ��ZG�c��z�q)m����C�9���P�0{T˘v�#�mQs��xO��x"��8�Jv�r���6�~�'�n���5�l�R�+׷O}���`� ?( ���#6���HT��A��$���~3iJ����of(Sh]�Pe�M�����dmZ&��+1!VR��{�>�W�����<K�^��d}�2��Y)F������e���F�>���^���G�97�0�<{xۦ����yC����w"P&
=�]���Kق��87�7h{�Spހ�B�m�����7Ʃε�ڑ[��\��ـ�;��eLgn�M�6�]��k��㌷��*s+��ޢ5��Z#��ePb�7��I_��ِ��/�a�΂;R�*?/j';3��l��c�b��]��#�Bə��\Q`�r�ivFm�.~]���>��@�l�H��&�������z!5��<U�q#iz>?j���eP�RȖ�g���6�h���3tP��8��SP�������&|==���?X�4p���'̋�Z���)� *[p'� ��xV��8f��]z��)!��t!�+�"�?�4"���WY�/�������z,�9f��q���gl���q�k$~��
��(�+<u5��uNAkN���%���G�<`8��l�=}��|�c�Y����e�i+�P�V�Fi�\�U1��6��A��'	�m�jyT+s�>	���6;���'��sݽ60"�T�G&}����W�wX��pa��Mb�a���B���>�qO ޗ��G�}�)`�3���8P'����*�AR#f����uq� �<�:����\��~��Љ��f*K0E����{ea�$(�D�E�e��尣;�.FQg=;W�J����tؖ���߶O���pSq����!����l�a"~��SV��:�U�&��.[��n۹�1a�l