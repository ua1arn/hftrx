��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga��ʊ�tl	]�1�f�ʫ���.�-
a���G�EMB� �4)��/��A�tA �aO��Nu
�	�d���,RaG�mkh���WE8F�k�H0���N���U�L�ܸ*`��k�VJ/��i+��	'߈�x�Y�lz<I���n-��%
@&��Ek�A�fB<���)'I2��P��"@�����b�b�T྽���%΢~��|�Z���i�?�����\#6E��<w�?_�1y�T_�*b��.��- �]S�)|��n�<=�L��4T�{������=}���ە��W��z��J���#���h�%�8�y|zm=�{#N�%���H�����`
������.Nc���~�}�'�T��t�Sډ��OV�2����W�F|v�p	�1�a��ھ�.E-��_���=f� {$u�K�q�,,H���A6�+'�n�4�� �$�^;��@l�o��PL٭-��AK��p~وϺN��-0 wM[��9��<U��B�^%%�%?248�>���t�����$����k��ӭFG"w��SV�gg��P�ɏ��yQ&�'2՟�,�h��j�ʀ$LkbO��cx��Qb��G{���Y�+�F6g���PV$���zǕ�@PPa<�N$fy�&(�8�b����J|�Z�0�t-�jAJ����=b	�n+e`��Dkuyىku0EI#���\��l7�>��ݸ���b��>�T-[g���@��1"���k��Ϝ���3L��X�U�?�Q,�)Q{h��U�-�B}�.�~�p_���R�ㆁ�?x	�B1��'Qk5P�͔W��CQ_0���L��y~T��0�X�r�ܚ���P��6��C��X\�i=�u�����+�Y��������WS��y�6��Z[i��Ero���ˍ���,� �.���6|}���A�!<$Ҩ�$��pY�=T�l���_�P�>4@r}3T�Th=�D$�:����k�����i�Y�/T�5�=d]XJk�����(Ub�[�Q�$�q��p���&DF��N���{F"��2��+[�=y,scn�V34�����'k��I�Q�R��~ojX�LJ�����Y�B<�_k@),m�_
�܏n��ۑ�l"0;S7�DC]���7fA+Y�]�Ô�~�k�>�|s:Yri�G��ֈB`&?����};�h�|�y��95aЏoL�;I�\G�HJ?���[o<�0G�̗P\.��I��w�y��ύ!��j�)Ao�S����o���c:�2� �ZXpv*L��/�5��M-�����3�(b%�7�N@ #]��b�*�eH����0��1^���	����6Ŵ�ޯ���!SP>�+���J>=�s�5b��N(G��Mo~�w���y_���Q�3(6z�v�k��Ҽi�b3,0Ln�����"n}���f@I�%o�Ρ_f@O��Hy��`�1�]2�K�se��˅@��M:��T6	�������r^ߺj��g��כ�KЪ9>�j���s�
u}K5Ih������h��VMW���K9[mc�����o<�ø��(,.$�{�b��Б�C� �cq�rh�GT�;Ͳr�i�1�� ��{��x��u@����#�Iӑ>4���}#�W��\�9��.v,��J��-oQ�����r][��H*}�L/��Q���}5��#yJ'�8��5���
��y�B�e���Z[�}�@Q3��v2m6�{tg����FU����,`m���(p�Z^!�8���7L����'���CXC$�Di%I�����D�X*�Z!�=u�F�L��Ejx0V���9�� �W��C�)`u<�]���p�}(�"��md��Us�+A/�0�H�G��J9=�����-�Ћ��7`���,%n׀����3}m���Ĺ(���m}Gux���{�X4Bl`Fg@H�:�;�uE	����m�O)Θ߀���쥫�\JYx����1�q���	����lxr3��sU]�����d��>$��{�P
������趝ַo�/;ϧ�!�D$hd��h_���]��ѵ��A+cP-q���q�Os�oo"�a���#z(A�(�̾�G�1k���A%6i�N����jF��V�*&㡳���V�*�9�o�M��hienH���q�ů ǳ[h�Z�~R�����	(�hn��/ 2Хm���@s�-YP�7����|3n\�o"Gu8����n]5�ag�|�������	�̰O��zE��5޹�ڠ��M��� s�8uy4	Z�#]���vo1��
�X�zZy�D��I�v�#5�/Ƴ���%6�<EX��PR7���n���=d��� M�	�����՞H�҈K��퉗��7@��Iյ�0bEUS���u�l
M�D�Ȓ�!�z#.��O�!�	�/��[��9MhbOP�|!׻O�E���MY%�C������T���]N(%�*�	�Nfo�5�]��q�X��٪<�^�L��:����nt�(�(��Z��t�;���y�B�C��T�����0�����]�a�{�z75�4�x�#��{T��)���S[�����^�Ff���_�g���jq�'�����v�o[��P���{�&��+���=����VN�;��D��$28z�>�M�����n�3!i(�����h���Y#W��J�Y��o���&^�T�(���mR
4O��q��m)�v���}�I��B��*�Ivp�� ?�p��}�3�5ݣZ�x�L˿��
37�D�8;ԟ�<����l�м�Z&�|vK�\ܧ�ˏ��f����0I�qd���֧)M-��I^��J�ä&���m�,��K�O�'�|�� �\6��Z���5��m�e\X���\'a�����K�*���| �e��7A�v����xy�6:M�V�E9�����^��A��p͆/K,�jEU���F>3���vUo'�u���?����� ������0B"A\�{��`Ҳ�x+�?Р�����i�k���H=���?��޴�Q�+Z�A	�S]YD"@<�3�KE
bef��
�;��S�)���Z f���W�"<�8�&��x�V�l����x���r�=�{�'�ԫ��^~2��XuЧ�K�!��0ś��F��)	��;�������>����K0����!P<��`�_�$��1�O;�-��E9���+v�����*O�Q�(Eק���Di���[�d��}��g�%��R�F��T�N���C� !}A����f�>j�Sfht%��[��P�����d"��ǟ$����W�ʗ#����W����σ��W6����P���WXd·EK�'����4�WS�;�؇Er�g!�'�R/�X�n)�>��f���#v_���� U�~[�f^����q~Z�}Aϱ7|q�Z����؆'�bL+
�U\5��dwisF�Vnv'tW����)$���K�j���w�����ޜz�h
'3%# ���;����-tڻ��F�ˊa���LG2I�2ô�5�����8�P{��ڌ��F{&.|��}&���,)��H-�ikA	9�3TW�uE~2�kP5��H��GV��)A}�~[u�U?ȯ�I���[�����a��#��H$!-ã�L㲃�9);;.5�|m���#��9�&��GSU0z�����M�P�kp���$~j5��K���%�����aVEm)���d��A�P'<�;��a͵xA��$(�3�2�Z�P{���g���#��`Kbk��Щ�Ղ��=[��t����e����$�"�JK�h`�1�p� ���`��א���&��-�V���m���/�fS�`��we��q��SE�q|��YVnO�9�wK�� 1|m<օS�a㳞V�=e&�mz$P����oj��YYJ���9���R@�n�������r�:b���/F�³���1���\G��@8��
)޳��H�{'ߚq ��nR(z��bpe�.�余Y��X��o��x��PG�'������p/�����W#�y��_��_�T�4ʾ&r��W`��e�5̓A"+���x��vWq�^4Y˓[���SU�Bp1��
�g����z�K�V]�����S;�7|W��a�k{�4��7VKlr��9mϚ$G^��vĀ�cl���v5lG�w��I��kcO�!o#�S����n�&���a� S��C}�HBʫ90SPl�֌�� w�"�8?}R������G��'S��?DE
�P�/�%Z��${ƷU�OG���/�O�S�,UҋJwm������$)x�[NZ�-z�n%]�Z�Ԛ�Ҹ*+3���F�.8O�N]	o�$����y�`b���ƨ[�S��g<#�\ӗ��ƫ�� ��
�A*S �ک�Jy&Y�O����j�1��c�L������`��"?�LAH�غ!��N7�Sn�u�)�C�CE/��ړ�G����[?�`��������h��p&	%3,d�u��m������[�ۈ��@m~�������{��]������r����q�mQ0��$*gz�%̨���Zk�2��iO��_���-;�.Qo\��ES&+������P������P4�N�%qP��Faf��ᵡ#�:��/�A��Z������������&L��=z�̈8�F���7�[��2��w�zV�����1�9b��&�]}���d{��q�`����#��>b���7\�2ݡ�msG��o��mD�Y�UlL��i6^�94��҆���bdS�z)�Mk8��¹��Q�q��UO�l��|<.|'h�4��_����EŞ=Z��S��Jh�{g��f�`�#X<�}�k?�9��� �ۃ
���+�<��Jr�c�a��/[u�Y?�(҃D�h+r��yB8}	됒��s$RSMp��.؇ϱy�Ѹ�*NV�y�a�c�j�"��z��r�}��V_�ƈ�3}�<-�`���(lݶ��j\�E�k��l�[g�-}�7�Y'��@����1Y�m�c�����C�A�l����Բ�N��NUrz�X�
�GM� �;�L��솼Xg�q�<c��&��U�X��� �wjr�}	n��sO �)>�*-��<��+8��	��F��G+V��	�u����!ѽ������l�+���t0ݓ�f;��4�q����=G�y�{��j�#���ח���s2�>#h�\�;�tϒ���A�En�_S�eo��8lA��ɴ���{�4�	J�H��l�_�%������_�2�bd�#{aj�t���\�͝��C ���^��du�E���· �1o �kͯPW��}	Y}��!�[cǟW�H�ԃ�Wr�.^g���t	$�d`��	q�C�j��P*�T��Y]��7K�47��/��8=GM����vo[�u�wG9�=#F�z̔p3{}�K���\f5bK���c��(�+J�	��,M�R`���z�oq,@�r�Bi#�Nb쨻Z"a�@=ˌ[H'})�\aUD�Ν���-�&���H;��R�(���I5R6Y���+�.��DC2�֎u��~����e��D������*݂�Pq��ħ������/^����ؔF6*���<�i���*9��pυ-�e��l[?s���ė]�5�|� H˼e�\��I�+6�����s���R(�o����~p���6��6R|��H5m�����RȜ��B��m]M�-B�f��o���7$�����N� �V$�s�,��c	�����/}�|Ze�>���t��=���ͷl;;/��Wh	�\U�G\�a�܉ڔγ��P��1��O�6�gȬ�{?�'N)��+/7w���-��^ONym��GV󊠹��c��Q�`�+,#����jP�����hS	(�U'��9t��+��]�cc�0O�NG��+���.gx��{⊿��|�Q���[+
�psu,�k����9��,���Z_�Bሆ<���^:�Y�%w�X;����va�(e٭��Y�m~5 (���v��� ���MA�RRZ�|d,��~���~���6xB9N�aU/%�LP�oJ�����bs���M��z��bJ��c-�����c�85I���mjK���_�
��BG7&."e�l��S7���n�M�N�e8��k�H�����=-��N��˸HYS���1\��r��xL#p���,4�g"��+= ϗ��,�?l[�D�#��Y�NW��dh-�2�fT�>�w��yL?c/V[�����H�;:�lڶ�Ml��`�u�;vEl�D=%��n�����\�r���F�t��y��q�&=b%H��`�n�D��>��E��}}�v�M�6d<dI%͊��ֈI[���Z��9I�JM��y��R�}��"cUWt�9�	�S!&ۂ���`�q+é_�{�g������7�v^�q��_��9���jm":@�c;;�������ؑ�����m�T^*C�L,�f�0������S4粌�_�{��C$<��WX�q��)��<t����T�u��ZO*�w�A��ۘ�Yǲ`���W(-�{�vߝ0�DF����X�����U1X���P[�L#[����&Ȃw�!=���اe��O�{=�z:{p�$�ѤMߨ�1��~,W��[11l繢�{�U���j�+�5��l:6ّx����!mtf˒������	���P1�q��x8t
�x9�����,�i��.C?J�>�o  )F?h<#���[�nR�m��fN=���	��O���6�n-,����(W�6l�=-����ܗ�g�vB�Z�	&����:ܤ}�$z)������̟*���x���l�̵,�W��0��./4C����T:��~Ξ���%���Kd�QnH���A)������G�1���?�k0sb�G�8�vjY.?�t���X���s	d�ρ~Cœ�>4伲<�%v#e"(iDu�w�Bq�y~��F�ޥ�����>����y|z�m����F/�w]�d���OW�/�z���r���Y�S��v��ow��%{+e��r��\��4s?AZ������G)�>�$H�F���9z[��|�ED�Y�Ɲ}��ө��X����c����x���c��)_��
�[�o�Y%�Q>�U�	^�W���-WN�DT?��J��/�Q~�@��SmI���T:uN8_�l��BÇ�/�j&0s���J�m�8��D�ý�G�ڝ�b��W.������)�^��U��	Qs9ۇ����
�T����W��V�-g}�)f@s�u�I~Zѓ"F
��Y���� H��m��z-ҽk$�N3�;C��%��7𫟃�d��z]�������8���c��YZ��{v�)�� �ҵ����o�[s��)V[�2�:�_�ڸ�����A3t&Axa�Q)��à�o:/�>/u���;Uv�<��o�H�w�'Q$2D���u�����*��Q"��+n�w�9|M���Tg Z�CL��1�#�}�v&�϶^g	��E�M�����_n5e@�GtO�@���;9}�/���>�J���y DV������e\/l�@6	�p��tZ���a ���6@�̜�*dM2�o����.��w���Yw���x	���½�J �;�Z/��^�V��q���l+����w�e#Ϲ�F����|]N�%<����n�����}��u�]3��jJ��c�ꨓ�"�[�)�	���(9"��'�P�r�4Uz��zB1��!�+S��t��*��g0���� ��E���q�Q\#|�tw�cfstj���҉o��T�}wi��$S��n�'��l$��)�bh@�Kȵ�\�7�n_�j�ht�^�{�iͥ��D�@��}j��-�Ac�9����;�UW=������Ex��]��DO��w��2�! �p�+�v�^��Ky�+�\�O�aA�X��ی��hEP)�6L[�L�L,���1D|�|/���.{�����2�ĝE�*>��o�~�$�izM�W�㹺��]@�����G#$�Dv���ކ@g�*?V�)�~�����l��Ȏ�{{2��������a%x�6{��o���j���#��O�+j��
�AcE�2F'	��8�FC�R|a:�kp���>o�[���;���[Fљ�&WY���}_��#����tH�����
�%"\H�1Il�rd�0�bឲ8�O_��I����2A��R�X܆o�ƿb�����!�Q
u�s	�R��l����L���W
a�A�x�B�pv��.ť��m2�]S��Z�������5�=R�ȱ'!�=���CT�%�7�H�h:����`YW�$w}�g�CX��{�V�C(�C=�F�H�Q$��6�&ۚ3� �$]>����g����2��2fU=��b�]��\��^*0�t|/)�潻Q��"P�˴��*hE8�3���Pv���S,�?�TQ�Z�Yղ��f��ڝ`y����&4u�	�6�m��Iwh/n��[j�������C�2g�@=���@�rٷ���E���Nl�jI�?�n!�
/�Ɲ~��XPa���~�mpf��Ű:�FjlвRx�,���)Y��,�j�c�2c�ݰqn?�+���/N�9�(�|�֢=�_��*N6��7��8���?G̭F#2�s���ngɒ�������f��Ȥ�]e����D��0�ZYu%oj�D��Q��V`�Zp��-�u>P�A4�}�O�X�5�+v�*�,�Ӳ�.��i�p&MNMS`��a|��]ۿn�d��M�ד%���H��t�I��/"@�ŝ8��`��>9�u���J� ��3<E����>�m-}mFx�;?V����*0I�5B��0�8,#�HB�|��VG�졩B�S��&|���g��/,5/a���ݭ����� �I���b?�����\N}�������)l:�̒t�Q�R�0s��E�T[���v�Y��Eo��ܮ����>{����B��쪺0a�+���g&��.J���]�2f���-��I���ᤷ��������'�Ku?<|u�h�Rݓ�f��{]E7:�j���C�d�����J�ǝ{��[�ǳlN�x�+g0�:�d"��H>�KIq�ob�N<���	�d�Sk��,{��ܜ�Q��u���F-����� ��QL�"�����	�Ci�:���|f3��?�n��ؒ�L���'��$�E�'�,<-ʫ�.�q���"=������0�`�����w#���9k��{������,\��� m�غ�Gz3k��眘�	/��!���yI{�Ef�?W%�,�����\�>FeCU�@xL���Mr5�� I '�6�&�l݉}l�w��T^���Nu��g�R���ƇAh�<p��KJ�ShΌLK�Sx���5�e��VdA�"�k#�3ZT��6O�J�,^s�ÄT`� nh3'9ؒ�
�[�5Q
��+�= C�\n���S�P
g�R}��+ӝ�GiF�TòA'#�F*]��M���
=��Q+������_�B�d��;c�i��J�ٗ��=�4�a*s$��.o�CQo�p��TV������No��/R�e���\�J>J��^WT\m6b7v��.��L'����Vx� ����/�ഐ���QY��@e�5��&��s,��َ�V�Du���b�箢��'�PyV�Ί�UG��r�tv��tth�G1�L�6jv��dd�Mg0ie������E�]=�2O�����C ]��b�]H�9j7����r�|j���ԗ����|��槢��)�&4ͺX��o�N5OΨ�`��%���i,�Q�����sA�Aׅ��4�-og93��y"�|
H※��t��ݓ.N	�j����8.M��{�u6��o�?Ua�'�~ AW��J�ч���	�tv$M��"
e����pj�kZ���)��:N��(6���x=lK��ɳ�J�4Z{_��ė�����,Y��h'>_V~��\g����q��A߆DQ�1qR̸��b4�=�~�/Z;&�8ktꝟ-���"�j���{�-��	G�W�u���a�/�0��«�ak//��.r��{����d|J�.n
r�4�Q����'*�I-���Ɗu�M��Y��oB3-qk@��PWc�+FQ���MOs�gkɊ�nߞߎ�O	�[�g6�e�ky�Әm�!�ܜ�<u^P򿈯q-�6���:~�Е���z���s�˯�\�BH��;@�6ޏ��HJ�<j��(oJU�|�>N�Nk1�y���n�SuS�16iY?�Ie�N�h�#��Ӵ�`gP-��[])��1�{���H�Wh#���N�\-���[bx����hmmu�]8�eU��J� ��s\,B��)�p���Ȯ;���_�#� ���U��c;�;]������Q�"{���/��[8���1|����V8���s`��ږ!�,P[H!�P#+� �5�V%U�`"��8V���x���
5�]	O0�%
_�6��lN>

3w4�
���'q*�=�"ӡ`�ٰ�$�4�e�����9Aqޙ�5Y���o��A%�](�"R��|Y�nN�[���Q~�U�[�����~݇���G�Qbዱ��������a�'S4�	�?��s"*��B�0Q�j��R޳�*�xkm1�FrR�d�̺@��Rq[2�#dv�7�oX�ޠ���sB�!c�V�����g7��W'-�����.�~vP�)kϜO�o�+Z/�ױ�8�;Ut�)�Y��X}���J��¾\&���S,H7AL�n��S_j�$i}�'�je�ppzYT>&,��d�|3�m�ͺ ܮr��J�X`�d��-®O l"��ĠF����כef�WP��PEr�d>CaA�:� ��>5��	������O`�D	Y���fz���wڿYSJaG<�R�]R�)�0����o�7��Q�s-T	���_����8�����Gd��^��gr+1����!�8c�UH��U��0�da��o�9Qi��<�~Ag�e�]�Ы�i�7���S[4��S�F �o&��P0� :�T����|�y~�5�X�@$�8�Nן�'!s{���bg���x�G=���UA�w�|��m�h�O|��s4�Я��ռ��O�F��<�wאs���A��o�oV2i~[�fB�'F�<"\�>�?��j��@�h!I��6�X���p����sS@�O�&6�NX�5�@ы6ݩ����&��YLwc4���I��H�}�3�eL不����ҘʁK�*��9i�[r��2��~�s��?�3C�x��FÒ>�F,���z��[s>���ߪL|���� D����F�}�� $&�+����z��|�� ��;���m\e��6\ģ�H� vC���y��xFgeF�m�ԏ�>����������M���j�d1׹!�&�O/���i�S��,��(7J^H;'��<s����	������1�����z$G�:��f`��Z$+H��X���)B������'gww�#��]��e��i��\� �ptٸ��n�b2��Ї��M�Q��[�����,L���mo�e�Vy6��{E��c�<��Iw;,x�eڇ;�Ԝ�wQ#�s-a��rx�YZ��_ꓖQ����z	r6�k�_�+@�&�H��Af{�g�yǨ��l#��M3�W��_�h�H�d3,ee�n�h�Q�J�2� ��m����U-�{��x�l�- ��˫�Ÿ=��8�C������2Ⴔ<��4<IvN�;I(=��^<
��N��� K)�Z�HR���J:�\�^����M�"�C;<�>��1�����󚵴��Ȟ��r-	�r/k�"��|��?��b��<Gp�"�!�pW�i���q�0�*5^�\�9x.� `mVQ蜸z?������D��O]7�����U0���y��߹dpǰ���䯕>�0��ne~B��Xa��$�~n����~ (���t���e�m�P���K��=��"�����@���:�q%m.g��>�	�녜/����a�����,b�ذ퉩`�����7��8�uy���" �M����&�,Ŋ��W �7}�qdo_T�L�����I�#(�Tz�A��<(3c�g:�p!�o�_�h㜞� ���H�?�d
�p�y�@,����W�oz�>���4S�Z���'�#������W-H��`��A����qXʈ��$8�椬	��Y,��d�[3M{+������\��(�M鬾���:l�qf��D�#�F���G3�������i %����:��
���Ȉ�`��̠ܖ���d���[-��G��ь_��@��nƙޠ�I�9jӍ>��*e>�K�j�@��4��ŀ�C���)?ۻ��!��5B�ķ�4���@u	��s��z@����d�S1���S��6�t,>=�Y�
"q'>�diÊ�����I�e��xK~8!���#���sk*i��C���`7g��ɫ��`�ĥ�)���V4���
+���`�r�`*��	Y4��#���Q�x^<�b2V}>S�*�8��ov�&@�Q���cZ;��:˓=�.�c&VBG-kl��`�k���Pkitӑ�^U"e;�f ^)�@�|��a��^C>�N�èA��6�r 6�?ў���.=�9K������[+�����QXG$�a����T���$^���ON����h�B�qW��D�7޺r��+���^�Ki�b��u�c&x�{���{vC���3�+k�k�A�	��!�$��X""ٓ��|�ݓ���p_e�������#��~0���V���� ����%+ǟ�\�nN�Z��`�Cw6ae�vCh��ز�ǂ��WT�xgB�ʦwz+��,I�5�x���=z��iӳt�+`��~"tgN�Ӈ</�Ȉyt���3�[��i��>Lx��!���"h����51��cZ��]x��H��#�k%Κ�UR6��h�Zg�OAh���\t����{������
�}H+�ʠ�l��sŘ(2ǘ�^��>Xy� �1�3�����v2dI!�/(M����t�6Y�S%X�'m<�wVbx��oλA/&�n��{[l�n4�3-	hR%�`v��Չؚ)/<��)cG[�fv�0��5Z 4#7?��Ҥ��Wʱ��`	,b�Y1eTV�$[��!F�|ˏ.�d�A��ZU���=�B/ v�ҳW��1�gfhQd�cv���S���P���θIgS�#3 X���5='F&p���M(��q��R)��.R=7Cj��Q,��a|XG�tŽ<P��LH,z&-���b����� ���@�7B>/qjcjf^�)������
]���6q�'�%�Y߉��JP&�=�'N1�?#;>{q�n��$.�rߓB�J�ð��&:a�-��k�Xa����޴�'J`V��p�p$Q`�����`�x?�&b��*{�3�̤ZI�p��̄b]p@?��}\a�n.Kf#� ��\V�-��dEV����'���%�[ȍ�p�BxV�^�rXV��=}���C| �_�1���/������d���l^�k�hC�%q$Qɵ������u�C��9��f
�l��m��S�ZAR*L����[{h�i1�Z�'2��I����'μ/��mh���c�e�Ь2T�\��)7�8g;��}|Ơ�N�y�;�ӓLVE���+x��?��H�(�c����SׂᲨ=b�D�<���,��nB��.U��M�^��7��d�<53�z?O$99�&�l��@Я���z�V�:����lVC������]���6ɅW!��6�k�Q);<��Q�ўs�����'�����_� J��`��|�]ù�c�#���^��$�em���*���8�l>�3n����]���<��3��w���P�;]�#0P�ܕ�������CYn��U�>�ӫ���.ҵ�c{���J� ^M�:NV�;ܨ��Fv�2���b)zO�a��Ӕ4�����ņ:��U@9 ,ݥ�-DC�#�W�Ύ"K&��/��T�֝��S�S�gD�I�,�tVvhWc���g�`Or��ݍ�@�H`	��`�X@Μ+φ�^�m�e��Ą!|����Th�P�n��!"m[�
�ql��9�R��yW�+21Dph}��;��e�>�6`S�nS~,�̅B���'��8R�b�𶐄|c���R���M ������԰��ˁX�?5G����w�Alp-�F2�_UO[�Hv�{����]r��/f��<w
��KXY��zJ�/�O',ԩX�����2��ۗKF�t��l����$Ee�KC���stY��iS*g��7=&cks�+�6��*
��dFRAx1�e4h)���Y�#.CKʅX�_�)A�픟3�ɍee���u�+m������z5�N��`*�a[��=�H�7u���S!�7��\$�*��Y�CN�S`A�8��n�a2�h�*`��(dp0�$�A����*�&�+����n�	wGgh#�lRB'�Al�v�P!�c���W��%�'{�n怚�t�y�� ��ѝ֙I�kFrR��.�M(��J��fz���Fi�i6�S��	Y�:.�]'KQ羕�{To `��!sZ\>�P��̳7�A����]�®n�;<���y�sD��SG��v�N@��+���=�m\[[�PNQ6S�-[(��R���Bo�`�i�ך�[P۱��9gU�К�Yy�;��C����_�2��4��SyV܇L���
�%�tu��+��D���8��n��3�O^�"5�����1�%�0*ui�_��S����Ԡ7���	�i�YAM��x��i�2������U�j�bJۏ�	ݲ�Mo�����Э���c_x�r���o���6g���?T��&$o�����]�b$�s�2WTI����0ʀ+x�p�+Z���wN�$�
����X�V&{���3��e9D���
2��)h|\��(6"������A�F��&�t�dɃLvi"6��\)�x G���x����*�#dc[��V�oY��C�,[.8�L,��$� ���Yį��D���`��zF�Ȗp��7\��
�F@�0=3[�/�k�_d�@�1��U�\m�B3���e_��(\o��6�{50!���C�yyz8	�W{��Oa��Jd2�"���6�z���P�_���m
���`�j0+��Y��'�rn���e��}Z���-3��\��$B�HY����wU��.��it�S��b��(��A,#���mx	��7����⢖�I}�D���e:�X���2��-����/�&�|l����*Ai�T�Q�v����J���щ�W��t�@��t쓒Qq�l(�m����ȸ�KY����-���y)�A��m �k����r��'m���W�t_�����c_>��(�s�l~�`�܍��{7y#]XL "�ş�Q'̣bⶼ�ե����0f�������t�i��'x� [f�<l�gz�7��˜՘ҏ��B$����%v�~B��hd�0~�Gw�Or(�B�c7̒���J"�5{9�V���zt<���q:)�S��!�	���n?��`G�^��{��MY)hF�����w`X����N�� nBo2�V�?�r��|";����,.��|b����e�)]?�����5*.��W���]� �.D�ps���"�8�-����M
�J�J�+�CЊi�@g
������*r��Z��Jh���_s����jgA�\!W�"Z�r`%y\������ Z�bq:�-�x�'8�(3��e	�Ds�-}pwZ�U���)0�w�c�[L�hַ�գ�~HY�ڸ��_3*&�.�pA��$�dZ����Y���)ت�qjz��9�/`�\3c��s��D�3�Y���O�Ը���y��Ǜy3�܅�x8��q3��lJp/�v�������k��Ye�`F�������W
A�v�'Q�"�;���M�_4N~�6x�. �T�. ��D���t?��(�}�=��+uxc���\FL`M��g���B��[}�ZDs�)M�9��Eƚ��A�����aXb���h�B8#`�*i0+�;r�摆��\�A�Ό-�K��Uۥ�����,�P@IGn�}gl3z�����Yx�^C���e��j�J$|�#�vl�4�n�&h��SUl[�𪪅k�9�
�}%,j��msH*��"����I��Y�+�;�w�t�p��W��ϯ��̼p��)�خ�5f&��x�I���N�E�=,�p�$AV���I�d ���`�o(�������a�^O�<Ev�ZV$|�؅�PV7���9��g��EX��ۆ���u��+�l�9������4�cXlz߄���^�N-���㗉{��O���:^٬�75�]�Ѐ�Y��CLtW��ZĶ#0N�Vpb� Lg�C��pV�$����ҥog�@������-�X���t��=���0M�?At�P���-:Ϯ��9��9(�Y�e������ X��An�Oe�]��}x
���w�����@5���7d�1���2���Ky;�$��䛉ď,��������?�$�(s~��F��}�������amӳ��� ���pNv��g��-�k;J�b)K���O�Vt~�;!�w�K��S���tPv��G�K��N���	������$F���'A��]xx�#�(_�����>�>�4����^�Bm���h�1�Qn�tm�\�V�a�
�O2L�M��(A�,��@�/�F^�-'7�A�p��`]��dw�\g%k�=�%T��w�o��a;P�-]�q[n�V���x����T����,֗�L��f�|(��
�,�y�a���M@(��FK7�!��ʴATl�T鶜r��ْ e{P�#N@�F5F<z�?���u������3̷S0�G�*���L�<h��=��jD��;��9J}�ta��R�����[���������}׆�W�F��������q޺���Ƹ��s�Žە,E��n+a�|f�--�h�_���/fo]H��xٜnI1�h<~��	Bԓ�ݝ�б>Myq=��j������S`n��4���/^Ɇ��p��r���G�ED!t����o���i��ŵqa3��|QKQ(�5 �Ժ�'���-�gp���y�n\��
�MP�E�MD��ڄ���|���P&�j�2cL,Y`�r#ڴڽ#��I����g�6�~6[�Zբ���:���o�Ԡ?��Ȃ�\�C�R$�!dk��0}j�=�/��Jw��Ͱ{0���X=����v �hP��y�����3�L>�ȴ�-��mE]nTQѷ�!����(>��Ds��-ƌ�|�����>d%*�z4�&�/�kՔ#�f���+�X#��*���ݑ�ni�(�G�RF��������'�Pt��տ��37�S��c</�6_�[���q�?sА���>C[ø���h5�2}�q�����8ML�z�t���I�Xڜ`an꤁�À���T��
���.�d�ݝ�
&�e��U��b� ϻ� ����"w��,����ٷ&y��!%`� Ir#�ȴ�b���4I����b�~i�R�D-��4�U�K�|�=��]�U��[G���n̅��ţ��;�sA[1 
ũ��Y���Q��^����&B�no��g)n&�g�EɟHn�������*!���sw3	�KY>��Ch��XTb˙��@�����!�#�r�7�7`�g_@�>e' �2����>Q`G������+TW��x_��K	�mN:�M%�$��^�m�Η�Kg�+�������.��_��X[�r��+jk�Ior���A���]���H������
[kWh��$\�,MC�R�=�&8�#��E�v�
P�����苻Gp��_빖*=��<�~kO�59p�p1�(�Eٿ�+�C�A6J�BK�:��Y�2&�4��Tb)u��%(x�P3?��I�Q)�R�q0�*ߥS��7�Im{��x}�	o����#�MZ�B��`��X��D�I�a��u"5k�Jm�:[��S�7�e��6����J�:��0y �:S��:��&(�qW��Y�dgSw;5y�uI�h���M��bW+�x�#u���9��t4�pɆxv�)�?��Fd�7���K�M_�F�����M翩`�	B�0?M�a�3|�`�o�O��Q�={p��e�����k�ZFx����K9�a�Ma���K��4�����Mx����$l��p_j�_Z�/������� <-MU�4S%��0ƬlK`#벧nD�1Q��Z�9)ζq�@��>��m
}�c��d��4�k-Ԩ�ض���粟�I���x)P.x
k���(z��ڡϢQ5����QĘA>,�5�_���G+�Yb���	����"��w���Bk�����Yc���mr�p��sr�oZv�~q˒�e��i�����9`苡;Q�)}~�o��j�M@���T$�lK�=#q_N7롵y���Bs�|�@���R3"e:P����L6ro`��2��-�?���-`������0�����wΟ���?QWyYM�"�|�!X>����N���q(����F4%!n-����g��\�[FܸvXI��XvZ�r���)J�c�A�N��N	�	1C�����H��A`{�� �������o$�?>�ddB!�,�o��m�l�-=������C���/��J�Mn�L��[�3�6��/��f���ө�y���˄���6OW��bC��	Zg��~e��c�� !�������4��� F!s}��b�j�Aךv̼��Ė}���4�Ձ�=m��L�UTEt�J�� r�.݆�.�q�4c^��p�
���Q��m��~���0O���� ��La@�s����PpJ�Z��e�����J%��%ݏJZ�&V�vze�`���Q9P��2��0C������:��Fotk91�P��ƃw1����Rc�h�<�2�d��Z>ၐ�L�}<��@��gь��WQ��D�7/�h/͒���m��8��L���2��'��|䀪�2.G�NNq
� kTV e�Т��!1�Pڑ!���m�H�
b�c�ؤ9��ˈ�N�p��zP�&��sd&;��d�aW>V�
�5"���AI?=;{2�S9h��a��J4�4�}�b#�#�T>0�_�;-<���?��](ڧZ*���˂5���e���$.��pjQ� D�^?��b�r�l��HK5s��
}����ӅJ��_�|�f�Ԕ���	����أ"�)AsOyH�(ڵ<'�`ݪ*`<�Ș�׎_����'��yऽ����9��r�)�J�	�q�IZm�Oo���a�à�G�D~7��'w�s���L�%�V��_z�ἢ�y������ߞ�?a�>�����T�b�H�� �􌣕��%��b{��:O��|���sS�$�Uu���ߚt������$ xm7�9a�j@��@.���b4}=�pq��ԉ�G[Z�><�C�,�P�Y�V�8yq$a���AIg�].���60۝b�(�a����?T:� Sxv���hu0�j]63�����d�u=[��j���_��H��UcH��qE��f�1c�1���Qz���O�^J�S�5~LE��Y.O�Ň@5�s��^�ҎD�[���r6ޗ'�Tz`�����Ԧ�cRʫ2�b��������kl@�,� �u�a�u2�Y�@ۮ����0Z�D�awBU_y������MKRE�i/=;-G�Ҕ�h�=F��60:=�b[@I��}1�Q:XcBC���w��,�{l������:l7~�n��d6�ٹ��u�R!�^e����eZ���?��4�FP��*oi\�`3	!$�8Zt4�Іi�=�zAC�y�F k�ρ�p�.y0C,���F)�/ʻ�so��P�!��^�\5syK7H`y6l�;�������0TMP-ݪ�E
�|����Թ�Yn�������3~e���/�wv��#�I�-����kyQ�;��S��ߑ�Af�b�㈰Փ�W�$|�q��wS-�(xL5X��f˾
��ri�#K/3b�Ymgf�P�iׂ�w�����,ЇdҤS�`݆�u3�W��ȳ$���l�OSƁ-��?ET�To�YD�N=�z��<���G�y~,Da���%rM +o�x�����0�X4��J�I�^R�$��Kd��������#�C�>��>KS�ےmڀvv����s=���%g�D�u�,*�x1��q�����R��l�Ch�]�K֫� �b��ع�-��E,���ףּ�n��ET�n�!��'���P)��Nj��V�.�͂�9s�Þ@$Mw���M��l�Ț���̓9y�l~���5q��U�G��C�tf��{/�/�k���^Ů�)�ɴ��q� V���>�����[�92z�V��2�'���J�օkX����P�70OX�.��ٱ��,b���U�x�\��!��q9�ݨϚ����Ҵ�����P�Y�_�'����%��F��pWt/ǖd�q���l���Ƌ�p��";~ �����9�_�5��l�h��w��yD���q�;}�k��y9�
X%��ӆ��WW��̹���V�q�U�%�HΨ�S-q3K���!�iL�3��u��(�OTP~�r�]O���&��10S�u~��m� �1V�� �k��;(����7���O��;�%��3q�6�b�k���"z�g��_t�t����!�1 ���E����58쓯Q,;�M���4{*�+}Rd5�_������ەz��]����jA�tr�5�!�ɰVYvQ:����S]��8r����I�B�q�ϲ���ѯpW^|��U�@6�����*�zVXa��,�g|S�ٴ���n~����<vf�$%���/*w ށÉ�	�_1�D��z&|ڇ-��{m�T����y&
��_�YDS�M��Mh� ����Lq��A��
]�ȃ�J�9x &�Y�8E��� �T�οP<GN,A��[G�ȣ�����y;v�5�a	������͖jhZ��n7�e������k6>q�H���P�R[W��y��Q<�B_�S�
CUmK���F|������R��F�t����:����뜼ʍ#��`��K�OPڊ]"�@V���q�*�l}����}K�טއ�z��Ă�E���W��mZ�:G^���5E�k�쬅� �th�]O�����t}�Pw�	�(JA�G[n�ע�_�Ȭ{�3�K��s8�B׆Y���<ZaS2���b�煿�$�$Y�Ȧ�5љ]+)�p��#�[�9X5"�����X	���*�����B�8oz��A����&�>j�-��z�m|�V�@�I��J�>˟��
<r`�?��/O��
lJ�I�P� �ɰ�p1b�X!� ��$M5��H�R�h�]��\U}w�BR[�s+��Z�uce�����k8���MMƃ�:�HV}r
|j�Z/��@� �Q<V2_g�;Q:Vg�	6͇�Q��$+���uC��u�����m6�u�y���a�dGn��H1q�Bw���֯�LQ��WU��O��Gtύ<b�mʄ⢃�e�S�nz/}�W/���_�'NAI�ܱWͰ_J3ժ۵�PO�R�꘸^, c����U�BA�q��ֺ���a�����Ch�����V$�i���Ж�������Q��7�V�'���?�1��D�����&m���AZv���>�bw�]��a��+13a���*�xk̓O;��d|�T�۬����/�1Pa�{0�DG����KV_�Y?��l�/��ꝫ̓P� YR�M�+KE�	)(ly� :X�t��S�⫭7�ёر	"漇���`�q[�¤�M ��z�Aa23Eeg4��}$����ـ}P���oJ�J� 2��6pd�5ck��7+�U&vWB�+��^܂?1�q���t����w�C�����]��ZX�t�QY�	G�3���A���o���!#d��!RJM�]¶�(�(�MSf�/d�(�d�mz��{��-y6��a��Bg��i�$%��fM���%��l&+ՙ��^�0�V��;3�vD�����NC�g�~�HO
����qT��L�["�:*��o�"Mڸ��ץ`��Op@���0���7��GY�_B�