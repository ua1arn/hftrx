��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	��E���u �
_iG"9���~��#?��F�1���P+0�>/�F����˕���'���I6܏��=�Bnw	4��6O����s��|�`=�Q�[Uc�	u	��l)��PVE�8���Q`s����kdk�e�H���n"�l��!D��
��*&>�QMn�n!������`d��_�I�4���,���vpɿ=�P2�$�Ą��Ø�ii�w+,�᯺o�w���Rt�ùJ�V�����ŔԶiȯ2�u�<Yw�O���dcf���������yC,?8�N�MX�u�~B���Л��	{��$�試���x0.����v�����cz��;�@̟]��.�%�Ƣ�wϞ�6��-����P��F��@����YLe�Y�x+�@p��E���K���� �	��F�h�n��	@����Q�a�وU蚼 ��u�����	��饛�����Z.���i�r��hu��*�r�Z�H��� q�6������fs�[q����m^b8����6I�(C:�����7�V����� df�)�#�b6A�� ��c�����x�@�ؽX�^q	�!5,���͜W5����-�u�93v�XڀD�EG�ki�qj[�K��Կ�`��5�����������y$@�BlE\�YPX���dd���	���ƥ��3x� `�N��� ��A��af�ҫ6�^����:[�ύ��4/7� ��1a�� ����_a�,TZ��@�2o�$3���R-F_���	���E���d��V���
e����"7nV�u�sؓ73��œ���"��ю����Ư��' *XE��+��Q���Elu�\m93KHZ��m�m�%�|�CR1��֓B��^L��A{,�Ig�G�~`۱&�:fe_U���v $�G�ԟ?��,uX�-yl��F[�4v��K�"+k��V���&�	q��Ad���B���-I�����Mi>g&m�8��/v�JB��1ؔW��1 �s�:���m����еje'?E��>&F ҃r�הo����y՞F�i�U� Qn��J4�ah�7k���8;�?�M�)I{�sj�e𜶢<9�QcU�!?<��	�F���Ó�n̽�Xה����˒:@�����疟QE�:6SCg6���	� vAm"*��M7[	��"�<�"�\�e��O=�r�{n�a�v���ɓRO�:	��$$�RMlU�rqV�Q]#qv饊;�(7�'o#E��z3)��g�W������H�/�9U~A�ζ
��	�U���S՞��;h"�S�J��� ��.{�`�|@�x�a�b��l�	T��Ka�����	����n�8/6@7׈�e{m�hpKe��5C�Ĵ��I�y�Y5b
��#���Yx�k�F�\�pKx�L��~���7�!�]E�݄sm�t����[.�B�)��Q��*\���}Gi����*��8P��<'͒L�gn��ᯑ��Gv�A{F!Bl��$g��9=H/p�k��}�l�qѴ�s0 ?m�D���?4*N������7k�X����V�[Cɿy���o��C�
��=���;�)�,�]�=�+7c�&}m���W �rR��;i����1���U����׽�׹���\���3�Z�J�j�o�7ዯ�l�*܊i��8P�J��U�j�+X\��/$�s���f����LhG�;N�BEwVԶ�3�p��rV�/�R��0���*S5��;�v}�I���~�/%f� J���<��~lp��}��,J(���k�蓴�k�Q�m�l��ks\�j��
ŏ��Ґ�Q�����et�}M�/��3^Ʀ^o�`p��WpNq����+
M�P�J&*�ZWvǍ&
�2k
�[s*8�8TEM����Q�1z���E��'M �r�ehٝS��6\����B�� ;�t�g[��~s��ji�g�x�=M0cj8 ��P/�  ����ߺHYIB�_e��T)>>!�I�c3Wϛ�}�`�b-��MJ׺�u=�/qC~��g���Zyޫ��QX\��)��&a�����)�zIT�s'h4:5Ty+k���:Ǉ�;w���o#���n�HvCeW+B[�D�DN_�hMK�~mצ\M(�8�? �`T��Up���m%F��\�fǌ��@���~H�R��!���Y;�I)Vlؚ��?��s�'4/���0j��G��}��K%zƵ�����k�H]�z�	��T��d���uL���o���=C��3C�,�a(JI� �*� e.��f��PP�δ0œZ{NE][Ŷ��1ڥ"3�����<y�́VD�앖�	S��8̾��oO�o�SU�澚���ޗ�/,�.د\2�dG%���6�)V�dx��ȁ_G�?��m5�33��̀��<f�!<�|=���B�Q:ɕ;M��,+�pr�lz=�5Dֱ�mg���a�Nڳ�.��bCO��=�t8{8��CWz~���^�C�(h���v>2�$y�?ڱ$�ˏ8��r�w�`�b͇���}6�� �]~�UX9N(�� ���DRN-<:3�%ӊN�X����4�|#s`���Kѹ\���|��pj�y�1p�KΊ�!à�m,J����vf��B��Z�9�>c
`�z��d��1��ָ=>s26IC��2ձ՘�̶~d�1I��?�%W���J��"4lx�� b�(}�m��{��s�.�YF?�\Wsb9�7,m��Q_U"�8(�!���a���x�� oi����:o�x�A�l�:�D� �|~�^x(����p}(��>�o�ucq�%9�vˉL
}l�.o�;�Yi�[�?��ɛ۶��r�+Qf�c�G���mP,�dab"['����c�����P�HnX���w�1�2�H�]"�~w�I�]'/'���!k\: O#��~�<��p� ��@�����")	 8�2oî3�Q2/�cF)o����]w��e�gOL���X�N~O�i���}:c�0̒�����������镞@
_,k���I�ěnyȪ� ]_��knLP�4bI����,@��
@�����Jﶨ`+�'Gy(�9�v@[,���0W{�|�
��IАqAN[Đ�m6�1i���Է28��G�ҍ���@=l6o�~#�ٵ7�Lg�<-{�7م�kl�'�����땰��T�g7~q�?N�������O.d�c��9��*	Y
nk]��Z��2� Ҍ=Z��H�ݭ��c�w��mhr��!���x5��M�,nd.j���X��������E!��؉�4Xl�k�u~�o�����ڽL$/|��\Z�!�������mY���]"�	�ܵ)��c�����s�.�(?>�7��6þZnN3����qQ�0K���qbh��td���6��}2��Ϫ��ω��]�qʶ>�����+�&�݆5ޣzk�i����DM <�q]�f�>�@Ɓ���nc�����dykz�S}��$�.��)��< ��!��x��䑃`qz^�X�#/<� �0(��&�{�R���!��57�$r�
X��0�d-�`��bIJ.��u�-Oy�	��83QJ�و-C��~�j�J����j� /�|4}B+@����g��h%Z�	�;^{>��]���IT��`�jq��KT�4}W�W���򫐫!P'8bٖT���[�ߡ&�{�Rx��7^<���#�{��"�>PEֶ���Y�<�Z1��XI�3U��WoW�b�4���ښ������3��p#o�W<�M9����;�pdci� �(����?Z��ef�_�I�J[�L�� ��}l7x�!��;��Fz���L&�n
�`c���i>+�1�;� N7D�R�c{b$T�ҫ�:ծr�SLԼ�| �F�֡�f��YI��S'C�I�s�=Tn���P�'C*)舎K�qUK.�ñ9m���Q�����8��,|h���9;�p	 lB��@P�@E@f@�˫)�E�:�?ɾ�(Ό��'g�l�/��� 4W_�����m�V?��G�%�,kd���G�Fg,�����KnO�l	'�J8�*�|J��t-JN_�6��x���?��442Kk�N*[�DN��5a$� ��bn�=/����j;\���(� �?/z$��ݕ��va�W�� ���8���{�/q��;ư&"[�Y.�%r��r�x!�uI&��T�ݘ打A�o��KAoy�@��#�.b���X	�"���9Ȁ��@��"�L���[���7:=�/�|OŐm�����v�E��͐n���W�*�����~npE�.Q��iQ!��iA��?���m��$�����.AK��ʛi�ޗ��:DC[��6R�寣?����Қ[��mi����0�P�E
I�y�c�yy��	������pt˼1�&�c��"@\`�������wt��O,gݍx�ݨWW��c�7���HZ�LW��K���T��`���şUs>=*����g�~4I�tExY�Nb��e���,3���v ����	��[]�(	 ��h$7��%(Uz�o+KH*�g'�Z��;��_����E.�|�B*
�6(%�q,�Z���- 5<��V�or�AJ�¬��E�
�~k!*�HC��z��29�W�Iy�҃x�\t�0���߮{�|��B@6�5�����ʠ�_��A�|x:ޓ��ݜ���s]�w�%�nN����x���y'�8�ǡrE��yv���I�%
��P��N�g<��Fg^9�5$s��Ό^z8&ǚR�������is��"TN?i9Ū��J�V,��I�یzw�k%�k�RB��%o�klu6��Gx<_V�6�qfn|�
����0����}�%�]��ۖה��ap�s��b��r�G��ɑy�aA�(���I*�� �v��i<��ߒD��l6\����mR}�n������$nnqd��kt8�H�ܙP���S���&�p�V�#�s�������t�.�3�8��z����4�>���脾v�������)���p�7��@�a��߼P�u~�.�������Փ��
#� �~ �1��,���;�)2:�k���P�ϋCPVrkjB���<2��H$�^WŒ��5k'x��;vzm���?�-B�؋	ìe��Yt�Dt����}�J�~�$g&���%���wYb�ИzˈƅkGz:f��J�������@\'н��Յԯ�&Ĺ!����R '/�۝��ϟ�u�2�������2M��j�q2�v0�1�3��
�@�s�I�>͟��?�n59p����I���ePF�ѨscF��r�	x^���`7 �/�8�S��0�/<uQ�i9�Q�>q� �_ j@A�M��K�p�H�x����%�����*	\m��|� A��;�{�G6���= ��Z���?�K��J��F�	��B&( zͱ5�)�����30��iHNsrR�k+�m�!i� K L(��C�^J��谓��7���?�;��#o�t��1��#?_�p�_-�a�wND�s�o&s��b��e��^A���>2SR�e�����=���~ֻҁ������
��3��M?�wq�1> ��,��I����d{^('�bO!�7J��J�G����Ͼ�3��[r=/������÷��_����r�`:�%�S�(s�� �ː=WO�(,Zg{�����	}~�b�P��(�&|l��'p����Y���Vh��P�K/����M��7v��=�JF^��z��g�R��gY6��(M�.����+ @��� ���-c�B9�(?33G�b8��ڤ�u�p0xR�������cwc��m�����
�%HPZ� ���CR�����$�)hbr��d) �Jm˙��*��:��+*��e�]�MR�L��|������#�!���B���Di%�G�z��u� �Ƅ�mT$ic���4�FR���!}�_/�zUF��?Ԯ�S����
�2I��cʭi�$"�?O�i��}<�u�WVR����k$�4a��64k�/����?���������ռ"A���0�(ſ^�w+Úc��D����@&�������owp�%ׁ��K��TN��HӠ6�݀��N��}��l1�IȨ�?�
V���k75�/E���n��/�4ױ
Տ��� ��4i�F�3dˀؕ���3���nX {a�|!;�*ff�i��_���3�����[7�_������)�l8AR�V��$�>�m�Y���`�_ʁg2;�y魇Y��ߕ���w�^@a��WC$�d���ӓ:��d��ױ������r�"C��j�/��u8~�*��"w`�����5����?�f�j�h�	�Z�v,�=�TҚ��(y�ϭy��	������[�������
�b�rf���_ǵ2s����&��N輣3����7�K�럴*P�lQ��f��������!�,ʦ�q��}-�Pn�А <{B�ϓ15���C�����葀�1���o},E屌s��rJ��X�2f5a���q��P ����G�Ukg����E���?}�������xU�p����-�~��(�<>�����vs]^��-Q���i�=+�,�xܼ8�(zT0�>���U|�|qI���l�IN�K'�kC�/�"F�lװ&7Uw����E��jd��%:J�{<�||���u�"���ڂ�����w����i���+	81^����A\��$wD��䘅_�Ŷ(A�A���.h)��@3L�.�$�a�2 ��ڏ�'�
���F/��QU��ȴcO��Lf�!�n�<4��9UD�����iRJ���"���%Ϝ����~+�I��qm���H �dX	�A�{FGl������
@�����JY%Jo�{�x"p.�[���q=����z�a����v�s���*Q�#&��)���SA�z��[�E��<�E��k1�������e�C�GN�]oHn��7CT@Es��GJoY�ێ��6;�u$4P��s��*%���*vĕ©��W����r�yu���O��UX�5�M\£Z�Kf&�y�u���6<�p�X;��V]�5��'U&s�5u�'N���S5��m/��\���U`��p�P�JR�q�$U')�<O�o ���H�Wj��A����O�QQ+�^�'rc)r;�:
�z@a�T[��w���R����Hʆ��*=���im��(����&0���,��n;�D%��s��`{p�_Z����\��G+7�ҩ=��4�\��f���&�FZ�1N��H�b;q�u���ymɉ���?R�W��p�x	6��c��jS	������fT�/8��.�^'��t�Y�f���:}�����d�R����g�a6yI\�Fd�9�Ė|�i���>C�]���'��Y۞������4W������z�gkSwP5�	7�A���߈�b��^z�E9�̜�B��\)�K5&ҟ <��Ф�/ԕO�vVy�V�ۍԃt�Z������K0���"8M��T7�����o�T�W����g�y
:Tݔ�����,;�~(�� �~�[��{;�#��}_�$���ֹ��?�� ׄ��LR[����|�x��,q��(�N�DT��%��6�
b������=�FY=�>#����N�z�~��D��tgH�MA�*�o��}�D\�H���6�0>��5��O��!2���o�(O��V\�j�+U%���)�$4l���z��o��w|��PX��_˄
�C���IG�d���bNx�q�o&��q��GdA2�mB�)s�I�%�V$�Q}E��X䜏$e�`g~�O-������k�Q&�C/+����*r0g\�.�����mN4�n4�EJ]Gh��ug��'�v�.Oar���#�� ~��,�2&����2���F�#��N?u@��~�;0[�f�!���mR�ߘG�Vp�ZZ��V�Qթ���Hȿ���3����R>�[��o�>]�uo#LJ��b�S�#��$�?��IX�3�<��!+����KVl��n��":Վ,s𻻨��S9�����U�ܻ7nn;]���B|�ÞS����]y�)?A��\�HC'�Rx'�����0���x�\�A>�h�
�>�K�Ye�d6�9�ln~�������A�ٵ�0 򴧨=�����s
?��u��L��Hʓϐ��ǜM�����~+։a"iT��"�b��c�L�}�n�܄�Q/i ��^?1�!趐 +"b�z�BG��6?��i�yIA0�<S�������	��(�� ?�|׃I�F�7���Y�7�gخ�ߦp�kdꩾ^�:y�!g�+lI���V9>�fR`�XWJ��b�X<ni����k_;� -��iqV��T����H
K#b�<�U%��H���5��&����T�S��*��=/��d��s�M����NR����	O�o�{./ �%�o�(���E+�-�C��~J����#�oJ����
���:}���&�.�H����9(m���8+�qg������Dv5R��ȥ��k�:���0OG�\�CX+�x�?�A��1��H�(L�|����qA<m޶L>g�}�޿�V��m��ܢ����.U���2@�O�V�43��RR�f10>��.�֧�f��_�� ⼇/��J�Ȩ9�$K���	9���Ϋ�G�G�,�Wj����D�p��#.w�jDiEA�o�٭m�~B!�"�Eu���h��Y+P�"��h��'&�Y$%4܌v.���d2s,�� @6It��׏���~�@qBH��V��� ?u�����3��(�q�ӑ�¨�P*�6#��#p���ҁ�[-\��m-�#�Sze5��z����x�#-�U��.M���,�jݵ(얾���S0�Y%~{�יwPo�П�p�[�a_�-�%�6m& �R�ץG��Ҭ���E/*�h 4�蝖>gX���O�JZ���,�p�Ê@L�ʝ: ��3��*k�?]�T��Eu;T�[�`ַF�
PP��q�ӮȔw�n^��'�[�q�u��t/�b�T]t�����nnr3����g��$����g���^.�Pڇ��	�k�D0sfN��k�y��B�],N $'���1���y�?&y|����F���D���CR�]�w�P|�EM�$)�1��	�h�����^Z:�>�����C������Wü��2e.7y�>��j�0|U���.ڏ� BA�_JG�L�Ǧh��L�аF�$��3g'y��@�Y`+���v�9�n����R|4I�b��K1�NL��Z-b��>�}�K��I����Is
�mD4p	�!�j)�"F6v�{��Y���F��װ0���U܆�7����\[0�g�"Qq����g�<ܤ�aˍ�g=1�[���6���/"��ܙ,+*�-g\!~R�.Hׇa�a��N�Y��~�$�w� �Q	l� �1޲'��ώ����U:Jp����d
��Hzz�7O��)Q�����4�+
 �N��-�m�q�뵀�8B����Y��)�dt�2~�px��+��,",���T�2� H�7a�+�CyB-\aU<=/�W��ā��!p^ɔcWi]]ER�£<� +2����[7��~����8��Ίp�9HÌf�Ρ��ǢkX����|3�A�0f����^:�xI�A�c��9�e�Y��0r(:�m�]�ϻc�/�m�a�O�[\���/80"��W�$�k�b,�H��2	)��>�Vls'��8;;k��ƶ�� fX7��� ��#Vʭ�j�c���5&H�e��T0/z4�?V��$D�I^����'^y��5U��zЌ�Mu�Ϻ��\$���ޤ�0�/���*뻅X�������=���>$�FߟRoʈ-$Ǖ����=���� 8�736�z~P_����_C��Dj�!��	����ˠ�DQ���,�a�c(*%�	r��V�
��Hf�ĵ�� |Ǽ��
.�!hz�[H,w�<Tm�A����?0��!��:��1�V�O�Yf��)j'M��i6m����B��1tݐL�ăs�/m��!�-�7�9�������0��{gVYh�(�t�m7T�C4�˶e-t��8�|U�m�,��b�:�g��'�t'�6�&�]�ek6��i\_uw�ԧ��#���*Ԧ�r���X	���� 6�r��� ���Q�xG�Ճ��_�9h�{tC����=>�������y�ʠLr��G'��[-���
i0u[K9Qt� #t�b�̱�,�;��P^�w �սڔ!3�)�  ���z�ǆ�[��l�&e��]
gꒇ��gc�$v`F��K�Ebo$+�E��B��Q�N3a�h�G��F�#�H�pbgGU"+ 8T�+�'��D����;�:]�um�Y�ퟣKq�	���:��E��ĝv�#���l��{�h=mԝ8)�Q���!f<��z�I�M3S�����U#��4�\�-%s^牘�`��u߄1>`��zg��PU�� +���j�����z�+�s�~}����2hAR5��2�<�����q�`�+5�S�N`?�;Vou��f�X�����"�,<�"A�,�r8��]tL?�TJ(�S�rJ���ᵚm�}�""f�p7���.�>���[�?]���To�����QXγl��^k
�)H���rXWB��W�_7��ɡ��H!	��;�Q���#�"��gxN)���0Y�>�_�l�}[�h�T�l�d��� ?�v ~v4���>/f���gʕ�g�6�;G�L������N�V�\�us0����uzY���E��"4㋝=�}3�ޢB���V7Y�JN˫Y^��Rώ�;,/$P�|l��e��zR6I����PL�CIO��z
���D�Q,��*X]�糞xɁ?Nͧ��q��D爡k_L��ͤ�	J�d�=m�C[�x��~<q�&�6˩�k�ɒ��sY��n�3�?����h�:>��&�m�E��T�������~��\L֬=֛PSjB-�S��{&,�ҋ�sT��0\ J�*o_cH�M�Z}E�#b�����0Q��P0a	6*��w[O��ߋ�ڭ;E4���;�9�b�j��aa�8lf+�ZәO�����ɩ��5��$T�Yu ���R��ض��c ��4I^��r"��4����[�gP85T�����5� �Ӱ&�I��/�����lW���:�}�h����+�3ɚֻ]��2|mqǥ`��� 9z�d�y�a}�-��{�l���"�� ��e��p�#�m½r�v����s% N��S�|�*��3�_8��fr{�aq�
��/8���m[+���Ù}��xoB�4�$�Bu??K:��,��촜�L���1�e�D#�� ������6?��L}C%^3����\3yH�	�Y^<D�9suډ͡yȗ��x.@$�@&Pt����l� ��᷆�ݣGu��RJ�[f}��a�`�n�sq�\u���ٔȶ��~��3Ug�S��{x��v�TT�9���g]��=��'��'�����N��<���	���]�z7:U�����1��go@�Z���|(J��Ւ�_PRi��#�qN-܈��b�Bt���+������<�)���)
�737��TG-'�9�Z$K,�������/��D�ܛ�P�Me�0���5^vE����*>�C�ǰ��%�p\cr�!OhEq6+T��g�����b��Mb��N.Qk�4��:B)����צȓ.	��l�okh�x�f�PADrʘ�*�Ob?�79*����%�U�F�wkQ%��W�*k��M�~[����--�j]�kJ�oM`�!�Shl��y�3��A��4�t �@��m@�z(�l/=�� �@���$f�h��/<�M^K�s�R�D��V���9hE ���n�r3��0Q1f�-�e���.�<���I(��4S�d�!<X�Go0����(�c�p�W#X���P1"r�?�>*(,�$������uz�o��<Y��%թ��0�K���~������q��y��g����я!���-��9�@�g�,2#�㚻ʋt\x�W�S��q�2}�W�B ��g�2��(3�I���f�s�N�]f@2�@�f�v��I��σ?E��y��4���w�%zҟN��ʓݓ�eO��_�e���ST���J�&�˦��@`[��52T�ӟ1�5A I�柽3�t�rSJ?��(�.l�>s�>Ja�-Q��x᥸d�߲Dt:JDXk�����v��K˰^��	r��\j�"F��{�	;F�������rAm�b_�fE~��{�֨!24�Oc�@?��D�Y��]��Z7��X�xS�a��];�9���n� T �pa���l�-ץ�D���>���-\ bW�ϋ���I/O��$wSF�abs����G���2v�?�6Gl*@���e�[x*�7��Fd�
���B�0��$�����Ǿ��_�d�f����s�:��H�0��,nh���T�ϋ 3lр�x�U��C��Ep1kj�Vj�k��@�XC����eT#���M�ͪ��jrw��bE��>�xs�P�=�]3�w\�%U
j5�MI�܃�,1�$�Qt�y��7=���o�|�GPW��!f[�4�2�*LcȈSw��"b��f�T�q�6rn�$����]�S��_� �hv
���|s�W�~< �_I9�������!np^gT3�;��b1�/��m^Sl˄�).!���B�5/gEKR�"�!��JF<6/�ӇEM����_E��[<��)�;�4�RO����O���j߂:���[�����{�[��F&l��<9��՛�;A��2���*��x�� �}*�}�yl�e
籄SW �����V�X��Y?1 ���:���"يo�!�#� 6��]D���`�FbR͍(����(H�|�e�!�*���X���%rDO����џ�m8r�Z�N
�s�/��b�+�&C��ʂSv���8">rO���n��d,
TK��A���=��T2���iѡ3�q��2+�qHT4Q����{�f8��,"��>���	
���Ի�{kW��یϊ�*���D���c���zn���9��^Ѓ�cL���N^��;�i��ʚc��8o��b�qg NB8���v"yǬz��E���"J��:O^�sh���c�J��"#��Т6�υ#F!�*��[�ƈƛ6�ޥ�_��U�(:.i���������/����\])�d2u.��0�	��uw���A�������R���,ʢ�>��h7�h1�"F��J���RζdTTZ�ƭRӏ�g��&@�Z��a%��'�^�~,GҲ��_9+���N�/�ا�Ȱ~xTI;s;U�}���0�pXF5ߢ=9D���|��$�+sz��ddt�Ӿ�f���O��mgV�������k���b��K�!�܀�l����U�b(�Y嵮�׫��n�.��c!���˦���-r�0��ub�1j�.�T$�BI�{������nL� �,����w\�q�"�e6[�.��w����k�1�hgaa�]�GU6lh�D�t�А�۔,iYJj�e�-�#W����XJ�7Q�`a$�����Hz]Țq�4�Qc�ݣc�&���*)��sx��8��'�Y�B�%���*K�ОR��|d�T�T%O6O~�]�^���хm�G�S|���+��8�c�Q%�,ng��$�d[fᐣJ�c
.���f�'��r�v|XQ����K�}���ys�a��@V�� ��z���tr��s.`*p��]�m�I��h��8#aH��[��]8&5��0�"�{:lW�V�dc�\t�û�"KMY�֛�|����"�u�N+Rj�L��X7�Ֆ(,�	O��6;Ue�{�Kbe��0�\G��_;wL�IIIx���ZFT�`���h��"���t���ў���!�BֺO�٧*ģ���lxӈ�e��`��W`X�~X��Y�U��)��5���=v�2n��k��/z2?���CD�2���;,������=zH���R�{�cã��Q��;24�हGȒݶ��DQ���N��H�RvQ�
0zq�����`#`u���!d��}z��+/��˶O<y���+?Ҷ��U�bI�^��!/�w�J�_� ��3��oŋ-��Vüu �1%��Й�|��X�)��n�3C=������<$FV�&,Q�:�NfU����+��-���'w���A���0��y����(�7%&��|B2w4����k*�% �Y��Q�LX�N����@WH7&}b:���yz���4P��;��a�R+�������l�i��j���[��2���as{p��uCVd�aҼQ��k��-�|�Rd�H6*���2��c�\(�Zs�_a�=�c��jM�lj�n$׭Ħ�*�YDi�OK��j�P,P��Έ��f&��o�E�u'��}/N��8��V��y��%�k/;oWd.ק3Q��FE�l˗��lH(w��X�{��F���6��d�2��w�����8��PZ��C2�Y��oY�q�`T���������!�yRg����'>���+���hXȞ���\G��/�I!�P�]YH>�<�ͯV��{3�[Ok:����\�}�mwXG\Q5}���B���(��s�*�F��A�S,�$x��/�O��SeJ���6�y¦A�Nj0��<�����:�WM��i����f��)�-��JqC+�_���2��`;���B0e��j�9(D+�UA
jz� ?+�Ľ�8� 'h��A%�5�fX ��^ �	��������.�����}K-25|��#�W��WS�ndG`q'�	5	a�$����;A�<ʰثiOtA�^�n(ݞ!M��KZwҗI�y4����f�V�j\Z��B�3򜎰	v}�>�q�,�q�4yOB6�a D�`�ʘ�g����n�l�2��N7���DOf3D+�;�9�0�%I��m+��$���o'��ȿ
)|3s������Ƣ��?�	�ӽ[��b�˨���L����� �_t�¹P��Vw�/;�U>��In0l��}���hk ēr��,b��$����l%�(��]��#1��YWGdЯ�S��(w��4{]o;MkT%<�IU�����P���w��X�F*���T�=�eJ�q�� .ϯ���0����˄�}q���I����N�X�V��Yб �i�΂S.��Rq��g0gLa2bx�e.�1�4[��N��00,0b��g�*��t#.���p�:1��Y,�:u��:<^U���k�:��eB'��6~�����FP�E�'��ѱ]&�A�>6���g���3�Y�$sqV`���3�Sh��2��y�Z!;���c��@����A�ƴT5��x���B>��P��(���W��I?	�Ec�#-�����A����
YI{��$���x��Љ��<�P�S�?�Ғ>	1V]q�D��٥d���,o .t���aL�-\�M$L.�$S͖�����P�_�	Uw��!l`@�?��Fe��V��r�9I�6�$�֭�c5Y1�Z%�-lF0�<��)1=>w��N)ܲo����-�_%���)���H��U'�0R��l�GU�0�S��l��g�d"WN)�1�����������%�z]�m���qϘ�ϲ�a��y	�/�y�h}���F��Z]����,H����D�u�N��;�㷳���QL�#'�=v�bNQj�}���V���9Jd�{a�o��vIʷT"������z]u��p�$]q�I�d��)��;�>�^��m]2Xۘ�Px(�F�>*�iEL�Y�0�+UO��h�1�b��H��\���Ux/���&�.���b�-M���ܻ�9�7p�R�^��S#a&
���R�@��+0��Թ2����6��i|	�ܼ�F���0��bz�N������^�Nޟ��"$��y�Rph�rs���%���a("�c��	}$M�"/�U��Js�B�BXW�õ�Ԥ���p�uu*ҵQ*�?���\,X숨�S����k�t��a���B���D�(q�c-�`Q�n��yd�������D��%��-�+���9U��(K�
��ж�bs�j�1������>A.��t�T�Đ[�X�pjp��k�z�f�������t6F���Qw����O`��)9�<�#�aL�l����!X�5�m����'BzhXHh��H��ZG�S�������r��}`ABư���lau��9�3��:~���(�mV���^余���9�Z�&l�ʟf���]0[T�TI7��(����(�xu&��X~�k�ꨁ{0���v;lSN�������T��zŲ��1�os�Ŗ!Q���l����e�S[a4 �.<q��-��Ձ�s��[����
��;�;S�=f

Z�u�4��Hbig6�������ii&ʾ���P1NDnZ�3":C~/����Dӷ�uXzi6�=-,��v<���F���d1%��ջ�R �ν���.�̡� �F�LZ:Z)��z��	
]wh��Ԋ�:�;��a
���=`,e�G�w3eQ�%���vn�Ѓ�V�P��ޣmq��3H-�n!�XɬdJ/�������}%�#z�X_����7g�>���
R�lv�+j�ف���W"а����<
���K���-�_��G6�ř��>a���[�XW��#�%@?�Z�����t!_�2�17E� ����c=�Yo�6�����3�]NW�����nbQ#��4E?�����(�}�% ]}���r>3��&�Z0�{�S�\\9�H4Q��u�|�I�O ��|T�e�s��D!@MK��@M�kmM���\ͬu2�F��1wv��<��v����t��":lR�˗Hd4�$`���p�� ������xkװ�"U�!�x<Hs��bU2U�}Om���=M{u}��%D.��f+H�J�
o��jv W�Gi����w�b��J���1�X�P�B��Fͅ:�=j��<�0�p�D�F�
UJ}����,��>a�<S��Һ�O*>�Vgum�%���?th����0�%�;2zz���h�T��i�Lbhf�hAQ�sUUٻ�λ��w�ꓲp���`@�'=G|�{�ǩk�RQ��h�zD)(i7D�svx�Āɩ󾙮m�nG�|�ܚc�6pe���1B ҇�>�2@�W�mh������P�e(�i�Zx�)�7����+�0p����*l����h,�)�F��+������O�V�D'�q,�o��`	��#���#�
��ЊK"4��(*XC,���+�� �tL.\3@��&�������f�H͍g�5>F��	B�U��G�>����,j�u&�V��	��6�s�ل��]u��=��7�IDz�������fY��b^aj�?�����p9�ܯ~@߂�R���P��s�5P�c-TZ������������?q��뮑=��_Ɵ�Ä㬬�Jm9�1���;�Y�R��Ы��\�roA�}7X�O7�{��<�����ُ .#}>�v���,v-T:����4�&��K1�O�j�m�	4�h��9�.�6��f&f׆�ࡡ=42�4O��>�+-Oʕ�d'�,�L�i|S���T��0ҭ�$�l���ǖ�<���`�L��MM�{�K,�0|�ĤSw�y?��4�W�����q{Y ��6k����
aA�sG s���H��Vn�bO���:�f��d�Օ���+3@|C9N�#N3M�4�ϻ��('��k�Zs�z����&Pm��� ."��Dj:=��ݿ��H2,�`�l�'#�#E�ic]_V��-t%�~��{���Iw��	W�+����8q|�ՑjU�:jm�ƶ)�Gg;��l7E�p	��xC�$���SCP�����H+���`��e�&���2fTp���F�w��n��rI�Ϛq	�� e�!�_A��4�R����Љ(���_��|E|�(��Ľܦ�y��yj|X�ާ.�g9o��f�8F�`����W��b������J�K�Lf�b��]�o�$���I���Q�m�.Q�E�ڒ��˛r�|��]`��!;���=X$c���+�}V>+Ñ�&|��%����~qP��=H���J!IH�lZ����#�C�:�"ضA�n3x�~aa�!նK�B0EI��[~�I>��B�(�xx� ���[�;�$ħJsl]��.?|�ĥ<��>'�����f���S*�>��O��t��j��I�FF���F��Ι�#���r򎘬��Y��-��"�Q�ͻs�{��8$p� Y/���`ҏ��T�L�i���R����ߐ ��}>�;�2U2����ޑ}�Pp�c�»(��:���`":� km1����حQwj	-`�O't��m[�F����F���v�F�@$�j23z��K�d�کv�7�&DL�V�&vCe=��_�\�wB� 7�O��'!�B,�o ��k����dW�!C���d���a;R�t�T=t�y�L3�&Zx�v��oK�"�0� �ӑ��/x��{~N���_г7�r=��Q����FO��a�����i񭎎���K�|�l�Lc���dR��1�Հ�2GIbށ�D��Q8�� `H��&�Ħ���d H4�f�렸��}ds�Y`WŸ�mФ��Ɂ�Y���v�|8����y���O���$b��vƷ��@8�ɨ¾4�i�7�}�g�P�����,L�^zK�h ��C�!�<A.�,Be�G�f�̕���\,�JL��sV�����i.��n��*|���P���ӌ�S@:�<akT�Re{h*R�M�n���ef�rCCAǪ<Wq�o�g���",q�՞6��9eAN�����	�ap��Jo:�=?
��zQ@��}9�FI�nkĨ7�L�&�%�B���Ҙ��Z�gтE�2)� ՚;�/�R��D��)�vdQ"�'�[�F�O���O"p��V��K�����^<z+��& �G��e�d�[�\�2�9�y��B?�0+`L�ȗz��1_�,�]*�z�C2�q�t��<�բ��s�����i.��+�O\9҈�h����L���-��5�Q�����Z\����Q'����,��Z}�9�=,jÂ��˘>��W�y��o���Y���0&�gW�ɨv<瀳��T�l7V�w�s(0��[i6
e��%��MR�6a/��K�..�N���1l����"���б�hp�mŒd�H�p�!M=��c0���$+Xqp�I�ʭ0� hJ4y����,�W�4�xQfռg�I;֘k^T�P�{��_�� �!aHdw&
����҂�f�O��z_j�qT����A�R�n?؈�!R��c<^&���0�.s��A��ɰn����
~b�'^ӫ�h N����+�2�(��~O�+�%��xM���K�i
����$Q��E��.���������g��v���)Rұ�n*MY�������C �k��/.(w�F�z��o��Ĕֻ��Z`�ES�%�X�]@�؁O@{B�X��D�Zq�_���]vu�GDUZ�$�z���.;un�S���:�bT�������3І���M�w�ʯ��b���3��4�2�mMK�����v��"塃�(�<ڈCzÑ�
��AՑEk����N�_�ҧ����v���p�t��@m���tO�v�#�a0�ł�_��Z�����pmx���a��@۷}v�}�2�9>LW1��u�lEy�����K�YnT�}9mZðr�-!�@�����!��S��(��~���s��͔�y�Z�[��3�KSH���+�M^i/�j�m0�KV1�:�'�J���pه�uX�)��Zf(.e%]�a%���#��4�����r�a� �!o�`��2���R��~�O�b���xo%^�U���4��~<T��k�eM��lO�c�dy���\m�4u�hJ$R_�!\,�PE�#�$4�v8h��K�@�)�6QIyS1�FQ��S9�Ir��׉S@�-��L��i�o@�4d��*��}٩]�/�H�!lD��&��˭�N�6~�6F#W/�+�vMb�.�MŎ��m�;h��.�=�W�2�$�;��X�i��,�����B��	I��*�Kԫ����AVU��l*�	���A�|[stN�<��C�7�k�lAM�]/#��Sn9���a�r��b�?��ǬIXv��?	b��RI[w�J��%UWɴ��e� F�g�&~,�L N���m�k�a��n����H�ʿ�vĜ��h�eV�r]w��q8@�={��a�Wd]~���/44!����<��v}��w%�BWڵR|��7U��ܵ�v�R)D߬�c,��g�#T �h�T��u�c��v��:�[7����9�s��3� X��ף��z�iGd,�d����P�7x>(��17p}��=22{<��1�]r���qt��ܙ�0�vnji%U[@�;Ц���m�-�2�r(W(.Hݘ^�wl�z��Ty��B������d}��bÂ<��khG+K�S
(����l� �a,��)����b�5�}��W�` ��!쇸Jr��!�0ē��ʃe�ԅ�_)�����g�Pޔh�br������=1��]�D^����}��+�S�����?���2G_�.PA@�i����jn|����)���bL�6�\m��Xb��ce�ln� c��,�%��tJ?�+�ڌ��ɖἈ�rPk�B^��ş���$��-oʇ��{^Tّ�e>dz���gu���<њ���ۨTĴ=t�ԓ����ч䠁�G!�5��]��`L�Ȇ���BBH_RWPt/|N^��V��pp��B�i�g���XIS����}+��i!�ƹ���ي�A�7��^�㙸�2�=��C�X������rt�$��f�Ȉ�R��:���X�vn���[d�-R��Yo�T%�
L���` x��[n#s�$v��$L�R�H��.�Y��m�R�ra8���@��sR� ��Za��F���)�L��N�QÍ���q-�L� 3N��E��]*D��}R]�$��b���39���YN�IE��}������N,����½��2�4�]�1�t�:d��B[_���<?lv	;���B��sPK�x�&��%u�d�5�V�w"]hd��.]��V�\>��/�Z�����,Z����`����j���4"8U�_�]�x]�.ܙV��]끴	T�o�!�ǵ�-,��Pr(>W���q�͕n��j&��UE����w�y�
f8"~l�Zm����:�pY$c��R���[�1P����׽�������E�>��w��wV�>��h�W>��L����GFN���,8������m�O�9���t��_)�H���4�1�K���0���--O\������l�ܻ���``2����Q(�Z��Q��2�D2}�A��fL\-.\�ѹ	��
�f0����h�[Me�����(�vƨԤ��ĈQlq25�G^L�p�M�q���r&ݐ�87��Z�URV	Q|,hĔ6��{B�U��C`���x����Ɛ���a����'^������l����楘Mb������e=f]�V.�a�bJ=�g����T�r����~59�o-7��@
ǸIԌTX��հ��4����A�H�Onま�՚�G�86&l�E�E�R�ʡ�C��{��j6��6'szl)�]h�r��
����`�:�%с��!���S�7S���]p��$�߰@ޗ�Y�3��L�]�d|��T�o��+*{�`v��q�����P󃈿����j8�0f:��(����X�Mf^�#�U�&�9�qN	漓��[���Г�����Nm����>�%1g\!Cp�i7�/�����e��0�I9���f�i��6�ڕ<��n�}�7�ww�p}KE|�N�TC���dsQb���M��V�qeK����d�&}d~Hn�������6�B��vr�<uV y��K���� +H���8}����ڗ�]X?��e�f�b� �D |�9ĢJx!����؈<�٣�(��s�}w=�vrȹ�ԃ��t'�{0 �3�Wd�
{�z��!�1�@b��&A�	����t@ȑ������$u�h��|q�`O��y��͜?�"�Z�s� ����,�SN�!(b4H^����"�m���alŵ'uM$���*i�*�/ݣܞDD�r�g����JO��XjC��M�#��>�3�x�1��j1 	T~'`�-|�eڝ�G��d$����dՓ-�5�E@)��u5d�|����h�v�w�������hm�h�c�(������~�Yl�����@ւf�KDI��D
O���q� %|���!c�Ja#���
W(���"�z��_��"h�Z:�ԗ�Q���3g6��H��)�L��I���3��B��#�8�Ŵo|s ��FK�?���ɥ)u{�͗Y�����@�96d���6/���(:$U�|r�Z����?}�V+�/>�=z凕�ڿ�)in����c{�ȏ%��+L��V'�m�C���;�ޠ1?ѝ� )�,�wj!F�7W�=q�XH��k�_؍&@9��M{rr��Q���Q3Qw��d�&&�%*Ң+5���9�]1�ͭ4���E��zD��DS��8'�����υ5H�_�F�r��D+q�����Mu�֪��)�]��0����-�^6@� 1n5�x�$�7]x)WCU������;�3?͜����{_�\m8��V��Ӟ<�CB���y�X��8�๰����6M�y���v����/Q�8�9�ϙ@����D�o˔c
�8���^b��G��'�gIU�q�`�=;1l"����B���2~��y��o%�u���j���/�3���/l������8 ������P����[�OV2:�{I_������gOC@�F��l;t����ؓ�?b�
�.~λ߃���zh��t] W��	�� �c^�9�-X\�^���%�; >&�u|Z ��G����ףO�w3fЈ����b�K=��d*rT��.;�Z�Q~����B����	�<~�pd��)�Eeb~�����w��%�T�����A����ţ֒�C`"W*��:�S�q%2QA�KO�HN�u���t��=���/v���V"����6P���s�I�7���\@hDht�O�Z(������c�� h�����N�!�-e̓5"�����&�O!3�9�����b}9��Ӛ���6qd0ZB���:�ͬ���8e;���*�auY�gA��٧^58�x%㐣�^@��ڀv_��T7)��C*��l:Ƌa���"]U�<u�@��v/
T������q��_��z��^�ke
����7���E��0G�;�m�q"^�)Ōu#;�.���N���^�$�l	,�]�KψK\Q|���X��� ���:��6}4��=�9#�����M��|'�"�,��=��3p�����+ѽ�hS�t��� �@�x������֑��
,2,��l�W�9���/�"��a.	���/��j~�K9�	�]�(i�ú6���?X̝<�_����b1�iC,�&Q�ڏ�/��30yd�˶�E��O�m��u��죍���֓dq-�$��{�^�^�sf�nR�����*%cP�};:�h�*_�����o��:�6�rŮkl���WV̈����z~�j��I�����6�%T3�:ϲ[7�D`�߆��d��Gt^J�8&x�t?��K����e|B\�'��$\P�a��ZQ�x���Μ��>�QOdiU����M�g��of�Dl#r��6TeFMXBCI�l��檩���*����u��M#n"Xz�N���@zO6pV|���DbgK:�]V)�?h����=Ez)n>�+Z��@�g�d���ܺ%%c�V�wU3�mJ5��B_r���^7�꙽2?���Ak��+V
��r�8�����5TKM�(&M׊o&ۏ���r*f�����l&�C�CTF�T,J��������X�zF䨯�!`�*ُ���{����Y��4t�@=�\��ˎ{>\3�n��B���G��St}}����������/�O�w9�C�,��`����'����~�7hDI5��������u(��B��MHB�I�샮BˍUd놽ٟ���i4�G�֫��FҧH=S��|l��f��0f1�V��uY��x-���pv�O�����"-��׸K�����QFI�t��Ʃ���_XHf�)��ɞAM`j6dӭ�>�)�CY9Z��6�d[zJ=�|2�He4�f�cc`���?��S��[!&xr5�!F�x�瀳'f���c�p�Z�m 9�~y��!�����աc%���'�.�3�U�y�_��XF��W��ә����xOv���H������YE��
�j��Pkf%�� ]R��Yu7u����q ] �����H�RϮ&�|���R�D7qk�g��EzxIK�,�Xi�!���NW89�^M��e6k�RG���WՇ��x.�m:ٿ�okQ���1|��Q����K<ƶ�{���i
H�=a����t��fW�Og���̀�bα�К%������X�r���4����{�}�5�z{,-�K�����/У��Q^�o0O!  z��F �ޅI�e�m�K����8,$j����q�D
���13=!�ۏ�|�	_o�T~��gT �����#��������*�P�����w5 t��z�`Y�:W�b)|�=�@��n"���A�cD�sª,��le^V@y�Q7�P\�� �;�8�\����H?Y�^�]:k*�qC�n�;*�T����	���nOs뚈���f\���$��RG�����c˶3��BZR��4�����K��M�������@w�������x�7�*�<��a�L��y�Fc.p�[
�k�\��6�U τ8��G��/��gb���<:���e�YZDCdU��>�-N���Q��KV������W��Vq�єf,��^��:*$���-pD����[_��֊�AQ��a�'��O�],�;2Z�^����y�uu�e���f=�i�8\9P��s��Al��tT��L�5D�B�xv���̐�y��M#m5(����9k�%�C��c�Ӓ����}0Z�t�y�|&�t�����h�>���y$�̡��-m5�����(_��s#�">�k=��Zr��2��x�Z���~�p���lR��.�����"[�"�W�UT�ٯ� �eBʹ}�n�=4G�4M{�/��ٻ���g�nV�S|���{���I#i<�ت���+ ����T�*����R�C�Z�\=Z�o=��i�^EkC�Z3�*�Wч^0/�YF�~d�I4���"D�da�Xe��jy�3oE	u�3��s��E7�r,���Њ�{3<#%r��;p�����gt�!�i/� �N�<27����?$f��>9�cJ�m�|�]�K�E;M���Mu0�)�=Q'���3���Ug��`L3��l����=?O���	X(�������J������ �h����IR!&O]��i�KAL=c3O�#��;%7V�8:j�d�}M辄�#W�j����U+��ͱ>�:�-��(�d��+���d��,�ߎv��V��42����-jR+߼�N(����#��X2�g�h��#���}7,,Zu)������d1rQ=��<B� *9�6���p�
�_������HTZ���xԖG�|T�*r�l�&��p!fI�0�!�E�]��%�=�T��0fh�؄���̣�1���y72�)���]Ȗ�C��hv��^�
���Y��*$�>f�v.0�7��2�m��(�p�?{r�:@����/���g�Rq���a�O��q�(����ʖ/�IM�uI�x��r�%8�0�/���o��:�[ٰ���I�����uP���qM�?��Uo6�q�x�8�!�Kh�ڒ3�3��n���/1�6�I'�`쀄�%�sk�H�����3i��Ė�Y�y�R�!��H.�p���5�.{�)�Cy�T!W+
�K݃����{���odp�н���'_� �ou��������> 'L��k��2Z�p-JV�]hR��6�ۖE�x��t����'�����q���B;�{��kX�7y8�G����Re]��g���|�V#bm���=i��WU�+k�cE]��ݎջO�k�\�PM�YZE!��Z!�h�ﰒv!q\��މQ�7A�I�\��*Մ�^� w�����Y��-x ����ǋ��s�}0�宜̄?�i�[���+h���@3�����0Qjx�!xʊ�w���\]B���v[��i5�/�Oݤs�����#c&�)K��u��>��A�GҜ.��cԲƜŨI��wU�-�Ch�Q�ء���>h#9Q[�,^�����t'W���U5���r�����U�<<��;ˆ���w��k:1���&��0�qA�-H&~c�/���C�gt�PQ]nkb��<�D}���n�􍠑>ZGx�@i�
2�q�	WO��?�Bf�e-�fk-1���Kc�V�	w��_b�&�Vɻ�| �5"��,�������ys0�5�))';�!5�� Wz��Ґt�BD/e��%Fa�b��$8Wbr�y÷�pˏ�]Ь�ի��	N:ݗf�)��w7�kW�#ݓj����ڽE�a��<�H������Q�#T��g�`�d#mc���Q�j�"���U,ʂ��! b�~�v��&*���l�����@����:�`<�I��œa%�_f��c�6m��Z����k HN6���Y�Ĥ��NAi�W�J����O���^���=��^�v���R������	&s�Wt�S������H/�#���D�3�~���+6hȉ��]\��8��@8~���W�U+�2
Haj�]�`U �$�ӣ�ʋw?�z��3k�����[��:���D�}3���̎Ԯ��s
g�$��O����ir(
�E]�@��"5��F���٧K�^~�Y<���$���)uY��EF��! [��N��)�s���2��뷁�ϒuP��05�Zw`!�r�_ƞZr`��iSm��a[d����z�=˹�
nD��2{Ҩ