-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_in 

-- ============================================================
-- File Name: adcin18lvds.vhd
-- Megafunction Name(s):
-- 			altiobuf_in
--
-- Simulation Library Files(s):
-- 			cycloneive
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altiobuf_in CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=18 USE_DIFFERENTIAL_MODE="TRUE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" datain datain_b dataout
--VERSION_BEGIN 13.1 cbx_altiobuf_in 2014:03:12:18:15:29:SJ cbx_mgl 2014:03:12:18:25:18:SJ cbx_stratixiii 2014:03:12:18:15:32:SJ cbx_stratixv 2014:03:12:18:15:32:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

--synthesis_resources = cycloneive_io_ibuf 18 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  adcin18lvds_iobuf_in_c2j IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (17 DOWNTO 0);
		 datain_b	:	IN  STD_LOGIC_VECTOR (17 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (17 DOWNTO 0)
	 ); 
 END adcin18lvds_iobuf_in_c2j;

 ARCHITECTURE RTL OF adcin18lvds_iobuf_in_c2j IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_ibufa_ibar	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 COMPONENT  cycloneive_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "Z";
		lpm_type	:	STRING := "cycloneive_io_ibuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_ibufa_o;
	wire_ibufa_i <= datain;
	wire_ibufa_ibar <= datain_b;
	loop0 : FOR i IN 0 TO 17 GENERATE 
	  ibufa :  cycloneive_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "true"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		ibar => wire_ibufa_ibar(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;

 END RTL; --adcin18lvds_iobuf_in_c2j
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY adcin18lvds IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
		datain_b		: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (17 DOWNTO 0)
	);
END adcin18lvds;


ARCHITECTURE RTL OF adcin18lvds IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (17 DOWNTO 0);



	COMPONENT adcin18lvds_iobuf_in_c2j
	PORT (
			datain	: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
			datain_b	: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (17 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(17 DOWNTO 0);

	adcin18lvds_iobuf_in_c2j_component : adcin18lvds_iobuf_in_c2j
	PORT MAP (
		datain => datain,
		datain_b => datain_b,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "18"
-- Retrieval info: CONSTANT: use_differential_mode STRING "TRUE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 18 0 INPUT NODEFVAL "datain[17..0]"
-- Retrieval info: USED_PORT: datain_b 0 0 18 0 INPUT NODEFVAL "datain_b[17..0]"
-- Retrieval info: USED_PORT: dataout 0 0 18 0 OUTPUT NODEFVAL "dataout[17..0]"
-- Retrieval info: CONNECT: @datain 0 0 18 0 datain 0 0 18 0
-- Retrieval info: CONNECT: @datain_b 0 0 18 0 datain_b 0 0 18 0
-- Retrieval info: CONNECT: dataout 0 0 18 0 @dataout 0 0 18 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL adcin18lvds.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adcin18lvds.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adcin18lvds.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adcin18lvds.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adcin18lvds_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
