��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}Cj�L��#]x�9�Ժ�-8w������G1n��� ��z9(�
jr�(-� 5O�`��K��P�=�GZ�L��#B����)��l��j$p�j{u9��7���R�qE�VfY�P�(�/ؚ�{
��.9��MҐ��9��WX'^z,,U3xo#����NN�0B�0�J���fh���dv
��(��m�ڵ�y��:�W�ZTD�)_ x������i��q�8*�O1�V�z�m���J��d�����_�T���?�
lF����O�����hi�Z�E�<r}��m����,5u\:�'L�[-���^��4��h�LA�����p��!Iyr�ipQ=A6����۫@���Q�/�m�o'�֋z�/1�c��\�C��NR��QX"�����C�ֆ
�.J���M��!�z5*;:�����, �i-@+v&R0oOGw���j���8v[��GoK�Z���^�\�K�,A�Z��CT����	"N� j�X�
�Y����&$4_�
�<�
ɤ��C]{m�ϭ=j���;��E!��2��`��ep���|��=��I���c���ْ�L�W�s�A�v!×�o�"[�'m� ��5��D��N~��!��U��/aw & ��@qjń�Koo���;��Y����+0��5���Bb	�!��������Z!���w�(�o�j��ܗ�@�fg��~�CF�3��$s������m�m�]�T������J�Z�~��ygc���睖��j�\a�q����~��>�R�����"�{�x�#D́Q�K�x��������Y���R�/l5_�i|/�0�ҵ7ͻ�q��������
�9�3s=
�`����v��g��

 #B�zV\�f��g�؏���t(_?Z65vQ�lT���g`�"�0���_
�����a!��"���d�n���򈰠�mr�l�|���������s��4�� z�����&��u��xF��7��5���|�Z��{���e�gN�Ȳu��1��}����8� 7Z;�kf9����ω�N(fw��?g�y�����4�^������']��ۢ���@��	��A��D�%�[0c+:�#v6W�VS�<��,�z��������Nx[ٻ�;-����z&:�b;ʰ��
@����T�M�dX�̖��q����������C ��>��Uߏ�[_]n��a�ژjk/��c'#Ȼ�(�!�<�sؖR�0�1/4����6E���������O�σ�w��I�g-�
�"y�)|x�H����;8���A��q������a���v�r���h�ǅ��tݨ|���Eq���P�s����8�`k��6<�/>ð���R"N���N�?��"�K�N�	�W���a@�G��v���|n����sa�Q���2�t�� �AKvt(	�#d��z0��t����ܘm�B ���QH1tp��,v�o��G�����h�Y�\l,&7!��J�+ϲ�)aźP t|�]�䖡�#EЁ��cE�A�&$�PTZw��;MU��7�tq�_���b�<�_�Y�� -Hk�'�"�/����5�_���פ��y��eH*��E^������3��&4a��F x�=@�mԲ-�����ƈ.*�������b*��9�[���/%]d	Dx;O�3ƼJ�63
�<��H)xU��1%�`��t�0A�S�uTQ	���e������;S�93�gu	�Yh;��D�f��8,�tѣ�4��Z*MV�)��Rny�y
,����Z������`1g�I����Ʋ��%T��Uғd-��nO����-�@�@�i@�E8*-��O$BV1iُ��HZ�*���5<�h&����eԵ��Ǟ��6�����Xx��F�� ���B֡_��	�< �,�x��B��F��5����/���Ip�k�����=!����&ךU�Mh��I �"���_��K��]$���l�Ɓ�
�@/ q�K��f���1H>){�[���d�Zl�&z���f0�Pf�d�f4��ʷ�����gz�+*��h�s*ſ���� �[F1���|����A�����~��09,�\�,�~�� �
�۝�[(m6��ǩ��0���YC�q���%�L���O�[�C��T�q�,ᇧ����$�A\N}K�,�k�$ld�<���]�%<��ҋ�QIC,n�[���0��&��BU\n���8[�����!Q�.��-�K�F`x�a`ԋwBj�EV
E�Y�&o��UM��0���-3�5eg�����r������b��z;0<ׁҌjz��>J� �y���t��e��*M��c�����m�ԭz�_���cH~AK�6|�e�|�!��M145i�7�",Ƌ���hH�9#��rY�#��Q��^p��M&��;�~��j#�Œ��f줲F<�O-�{>�àQYh[�\r��C��/�UZ�T4#���E蠸�;��.K��s�3� !�y/���`��s �-�a���3	�xX�g�*���m���z�W���q��K��A1���ܜ.���vpv&f�S>��'��uu̺�-�Q����W'��Cr��[.��֖����O
�&qgY�{�^ѥ�?��k�����W��.hX��n��eҲ(b��,����l*����� �	fd�S�!���8 �Į����#j;�G��*٣Z�fs�җ#v ,�����A6�җ�Ȗ��}N4�������3�'����q��iֆ�Lz��{�5\�w�J�U���P&�;����*�j�7J��=H]4��h �"�0#�j!a7���nW*{г�x*�ɵs��`iU�t��h����tG�&�c���`��+�_٬=���N�J�HF���$=z|HK���S0�I�=eZLsJ��T�׃�}j�Mh��c�����1!z6/������NQ /j1���5m*��6�GM�0��g-�l�-��P%BD�&���S�V�X`V6G�`3�U	�/jtT��ʑr��	<��a[�fW{
?����h�z8�P
s#9�m�{�]��j6�̀Fs��H|�nd}))��,�EQ��"�(Z��-�L�Xf"��{ڥxϘ�v�&^��?J�=�W��h��>�ucڷ4y�}���U���[u�H��UM\��d��I�l���c��h���˸����1�P�]��MK��6_���pQW��H��y���
�\�R�����iw��-`��t���No��"���iyg�JT��N��=�|O[�f~��)�lZ���|�6��>0�(��� ��c�dn����Pv������o�&�|?a1��pD�/>'�/I�Qz�\�yw�Z!�i�3ؒB6��C�J�^�3�1��_@Eu�Tsj��Ďk�ǩ0Vl����K�K��]���C0��5h����2�'a�9���-*� %��Nm�Э��9}я�̕XT����55wP�;���^�������Y�e�Q�a�Xe~��Xj��V�le:S��:5`ۊ�}	cS=>]9e`�Wql\ߝ	A����:ݭ��tZ��?�P]=[�U2�a�!��)�,˃����z:
�O{��ƘR��-Z$Un��p>��e�b`��^�!&��Cx�&ll�f�H4H^�����z��KY�ߝE[�ѐ��>�i=���}��Sij��O5�:����+�{�O���U=Z*HmE��S�ht��̻:ˮ��yH��̎XuVR�Q��]��C�⃞Qj'8,I�ܖ���la���F�4�������q!���>�pA|��+�"փ�Ƃ
ː���,11��\3��)�N�[G���N%�:ڨ�����^G�3 ������)6�'�/n�5J���\�@K��Z��Q�'^dsN$�=�Ă�z���b�:Hr��)���<���ph0��V�3����;!ǃ�����m���C��×�E���M�}m�p:��N�8\�e8[��r�u@7�(%$���5�J��1�[�礷*�(A� ����]���[���k�sg��*zL�ri�������� ���2V����-�;	lA :��R;޹&�����6�O�g�c�qӪ.o^�ڐS'ўyxe�7�l2�p��X������T�*����"�L�%0��t��+�GR��J(.d�('rZQ��}�*���#c/�`x�'�ʮʥ�EG@����'e3;�h���逾T���d@�c��*:\�����TD��P�F ��>��3����M+c��!&Du�P���P"w�E��Nr�8���v��],ɍ@;�������>��ϋ䓰���ggߍV��8sE�~��k�����G<����\�BRJ������l8��M��7՘x�X�=A=�������i�e{��e�./��l) S/=��<�3a�n
��l�����W�M����[��[��O��`�!�,q�6�Ǎ������	�"��2���x�EZQዸ�V� {O01�1����4$<0H��@�#C��VA1���"i�E/�����Cسa^����yu��W�脛NW[<%9k̷��F�t�Yo�/B�ª�ܵ��"�b�';B���&SUhDI����*���=�H�ƣ�q}uY�((�^��>�23�Rt���Ћ
��+�6��u�0F_�|��5x�~i�H�2	)�?�-Nn���/0uI��gd�UE"K3]��@�4��>I ǨE�O�N�L���Ou�?N�I��8IQ���ܝq�Kr������|(<y���P���D�� g�*7�%$oİt4R�N#��w]�'�Č>)��T�t՝�>����u�������R�F��z���+`R-5�U���u��t��/�5���G��+�[V��ޝ��p��n�~���]���>���t8���W���##�.w/�0Ii��M����p�LsU�Ω
��Zh0c �  ��1j���y��#I��sHWT �Wɧ����D�v�fE���[Mj_��q�$M���_��*�ⵍ �#C}J�e{����E������+]��҈4�ϻ�r��]S�f��ä�����d��F�i�D�hH�s!�S�:W��a
��Ľ������^�9�g�;ltgN_�*h�V�Y�޸pV�f@g\���]�(�8�	O��;�	M��l��Ƃ����خ�I�a��S4an����4U�v�T_b����v
�CT}n�6���e��A�ں�qIT֜��Ne�5��@��ޏ��biV�y�Ԥ�7�gI�]��<��5[�}����2���W��"|��.��G�N��:ꝭ�C�{��MK�q���=�:�Mvm?�@m:a���z��^	�exR�T`����!���K�:��pȖ�.k���T䀝��z�c,��5�"���vW4@�ۇH$+ *g�\ך���J����.Ŵ��z��7���\��蕃�����Q�������$�������G�A@��ȥG�*�`���D����2M.��շ2����ln�ñ��o�(Bl�@>*��cs�/�o�˄�d[��6��437-a5�	2 �F_���(�,t��*9������b�2�E?������:å�Bh(�9F�B㰹�f5pq(#ؿ��粊n��(	8�%�J& ���3oE���	�Q�B�9c��2]��@���l'�	�����ҝ�Z��\�h�~��H�9�5I��˷9BP�'����fB���iD҄|�µTR}�����RQ!��7+Dg�uE�H#�s�c��˼rϸ�+Us��#d7N��~x��́�&4��w�DOfuZ2��j0����m�s��������a\����.����kƕ&PB�ѧr�~�����˶=G�½/yeS�;a��NF	�U��1ھ
ҢP��l��Q���\�6�-`�
>������X^��P�㽏7�I��h5C�I��K�ܧhs߄h��ǹ�K9��U頡��b8f��N�jg�S����Ҝh��ܪ�$�O�db�dJ��n&��#��Q�t��'�$����~���:a�Z�n�z�E��Gy���Z�ϦY��|퀂q��jdP7Mv��Z���5�ZS-�� y7��ۯf
�v��a�Eq��g�
;��q��P���&�V�} =X�
�Y4����P�|����/��#�ha�03E;��a[�O�l����V�>-�WTA���ꗣ	��6x ����3�?�m�on�JtU���ǮɋJ�Ch�=t�#��}��s2���=��Z�*��<�ג:5DY�r���1>&���8����v�c#ū�{|�>�w����ȗ�&�jF���q�$�N�Z+9�?^k�v
Ǝ�:��Fon	y��fNՏ�|s��
��"�q�� ��T��3JJm5kc�p��H�>�)�	������E�+����%�jk���3+iC[��MH��"j5 ���s����v�7�i,1i���*o?����4���Ȃ�u���L�j�����3@#zU]U���@��&Fw�Q�;,�a����4䤘�L1!�5�_c[�+� ��Ԣ�����tB��5W5�T)�	��������C.<�x���"�R^�m�s��M��8������E���ˀ�X�S;�����O���6�������eP�Z���Mi�k$Z/�bo<7P�lOI]��QK`,����5��f��#�
��}З_�,��	K1)%��8�'�X���oL\@d_e2��q�r
H�Gfo�o�|����p.i���[Ў�jo�}�ǀ<?FތOɞ��w98�&ROtRr�˷����|��j����z�ǒ���QA,�C�����Gn1Zt�$o��#r��}+�r�6�ĭ`L5k�F��f,5�[7���)�eҖB�i��<Qb��ɸ=����fOm[��.��c_Q��� �<��e�~�`o�6"(C�5���h�D/ρf���q�LO�X8��+b~�zo�p@�S���1�6G��>���~+4p�����r�U`�ؓ��Q?;ks�s��凴��[&	|A�O�%����D5|T����Ń���v;��V�@���5�s����=�k�t׹��9�U�՜�:�8^��7���BD[a�=:��O�u������ȸk户~8��#//����0"�	�����CVJPz̮��2������ǹ�_����i�Kہ�d�t8�|Ūi�_H�I���;�C�*���vd^\y}�Z%\�`�Ҝ{�W�m��:��{/p�Ck���w�����e1�Y����L���{�^� W�p�1�c���(���ӄ|[��6�T� �����p�vlj˚���䦩v��/�_���!�r���7 ��y�z+��Լʙ��W��c�����ɷB�f����i�i5�ՉO�f��' ���,�Dj]N5�!�-!n�٬��M�;�?Z�^����Ar2��c�cG���CPv�,��-@Ѹ���ǵ��R	��/�
�5$P�DiN�2*��~5�â޸��ɖ?O\���%.f��תӦ3~��6���Ÿ�K���ur�8p�~�.�6�.��?��\�s���C�嫐���A�)���u�A-
-5�񍌏�+Ysym��rzR��
�]f���Vks`�!#7m(��r��+`�-7��w���ww8�Zu/$n��ZQ���Yt~�U蓗G�t_�����|�ޏ��Vv�Z惷5�h�{s������w⊴d_��&|x4}��]8��gd/7l��Up��ӱmV��_�౨~|���@������!��*��׍	M����p��0��)y�c�>����o��̅�)�6JV��@�)�����V��T�}\���d�\+�����Dk5�:*��R�Ur���LQ�>���_:�C���wR�qz��;ާ�<9�����R8����%��#�KƄ`�p'�<���p�q^��O4�u�]��ό+Et�F
�Tr:����|�g�J�N�U�q���1Ԁ�,-�LX�a �Od�)�*>����:��(B)UOUg<��Y�gQERe�"���O�A�'��p�/�;\�@D����0O�����&��o7�r]oO ��R�!�m���S�<Ijho��2���C)�Yb4���~H!�}f��2�Q�$A(��M<��4��v<�t��v+m��h�O��N���39<꺪;���"�5��'{�'`!����� ��g%�J��{ҍz�.�(���QUxvk��@����:U��nBSE�R���ݛ5i5j2���[�I tѬ��R׊��Vg�X�*M�����E��I�[4I���r(YM�"��'���Q� �R�g��`oLpC�/r6�&�k��^��O���4���g�l�%t��p@�i���A޺7�h}YvC�ڒ�.��`%����9-��+2�"��� e�_^A�A�d�7�2�u�u�(ʣ6A�;	S�٠���#���Y��g��>���1�޲uz��p�*�_LR�$�&���Ҝ4�m,��F/�,�T�	��2@j��M]���Κ5H�@�����G����L�s�F6���u�f�x�w�鲭��p�% ����gz��	���й���U�a��Q��۸ީ:y�FU ��Ȧ/4��؀OYLL`:D�Mjz)[�iz�O��k������r�ϾU�!���pP�i��%����=n
�I��v�htH����4�m3�|�HY���5��RP�@���[}>��2��VQ���&<^q*�/Q|6�ր�+�$�q3:�x	[���8��u"��j��wnWr�ʁk���|�ũ��hӦP7+n <�ظ�}��&tJ�qfھ8�L�SO��3���"wU�iW̛*d����@/������j��1+�`�q�ը�);�7���F$�\���R��0��=�XAT���Yf�=�μ2R���s�k;��>\+-�`�&��D4�Qt��Mkb�qw́��_	�>��>�u�ҏ�x��P;fq����k=!.BJ��a6������N���Ҹ��y��{���q;+?�e�f���7��hڠ�\:w����L���O�O�]�fBS*w���=8��F�O�Z�g
@�Ff,u����G' ���3t���G�;���`�'�G#�z�}����w[q���k��'�?k�;�ZH~
s�tB�Gh	�r?�� ��47�/�n�lv�bfy�V$f�v���y{����3!`���K�]���$���ѐ���(�1�$��;��U�&�E���������:���m�hfr��<nd���}7��s��[��������"O�*�cj޴W�1�&���Pڪ��̪Z���C�L��hh"�7��q��fv[�ЁtuJGotg&�`Rʧ�^��,Y��r*D�w8 ��(�T�԰�x����s��CΦ���w);LK,[�zH!��A���H��#��6sl�K���v݁;����ɜ���4�J�?+>D�-�d���692��?�: �$�	o ��I?օ~�vʃpm~�Q�/ً� R��zZx�{����륨{�dl�o�H
Z�;�jFIٽ�UW�)���ZIt*�)�i�e�� TUp�Q_v�,*� %z�N��h^���0��Qx�wb��L�U�@#q6)56 4��U��p5�t,�C1�&H�Bb�٭��p7������l�;[-��9�6?we�.9���_+��ʒ*��<?��t��r(t/��60牷n��F}6�~�2I�6.��K�'��%��N�yc�	#qպX��) 5�*��[�B���L��M�"�9��l��	�<^?�ZZ���׹�|il�J7ꑋjPH��x���)0E��_{%o~�jW�.���_�/���y8�u��߹�Sw	��I����� �ڳS�3X�"���BfO�e&�ak?�
U �o�2gJ�K�Y�L�=ںZ�L����X�����A�D���N��~!J~f	�m�ARy�7����cA��ڰy�o���K�Q�>\s@��3�GXq��\o���,�^_S�]n������b,U���F�(�S�Loa�»R�v��3�q��'�������pJ�Bm�C�kAn���PP� c�Y�l#�B`�Ww:�����[�������6���%�c7��K?�\0:��%�Aa�]i�j�w�_�D�}�Z����x&n
j�lF1�Z��Ӫ��嚌� R���ruA��FB�7{���󞗴y� )B�-�k����n|��u��}t��)E�SR�@�!�W�KI�1����:���lY{2r��W �F>���S{u�����sW'd���A�Gڣ�%sD��Gg�ǭ�D����u�*n�뒖��JJe=���eE3̲��>z��"��R ��h�r��0Y����=�,N�!+�D-'�s�� �+�bS
�i��6�@��#^R�j\0G^�Y�!r��S��l�����Zs4��P��bÊ�X�&�o�����;O���MɆ�\��%��!�U?5�k�̄��"2`�g�i�	*�t3�w
�x��$E0nΓ�E�����u�����lZ�K�A��6?��mx/R���l[ ��Vc�j�vi��o��=�/�����������="7��`+��F�"��/uw�S�Qީ�w�w�v���]�kٸ
F='�C2G��2R����μ]�V��W���{Lo�J4����gw)a�-��L��K�vf��r/V�~�f-����(߻����E&���>?���kj{{]\0��\6�ǜ�8o��Oy�.F�نP����r.6,�j�&��g �*~�F࿬��\m�u�����yr���_i����+��>�	�&�"�3)6��l�7km�x���)aU����)v��yDSyւ���w��G�k��^9�����ztL��G(0Αf�7��i4����5l�̍8����3�L�5�M����d�V���I���ӹ�Y�"����p�7�Z�)��ʎȦ"��>��|}������ڛ����Vc�2~N:�|Mt���5�