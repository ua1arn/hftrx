��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�X�C�[��"s�و����E��d Q��Ϝ�a�6+_�BC���~�;16F眵��bW.[�֤��%5�yY�v�U��/�h�*����m�0�5{Bǜ=��f�����~��2۟Yy�[�xQ5��-�Yi�q��;0|#�i���U*�{��~��z�� ��h7�\b��;g�aUU�s�����)�MPL�Ӄ��#�A(��i*�A�r_7�k_w$� kI��T��������Ul�I�-ۺb����inO���ORn*~Y4e_Ƒ
��I �7���DEt&O�o����Ϊ.��If��"�$�a^�L���|�$���o�����3���}*`������Hb����mcԆo��\}2� t��������N�+�U�r����5I֜�3��ӟU$�b���Apb*�����G~
��S6�л�E�y�S��u7�!Ȩ��hi)WX;&����^G��32����D��bJ�/f	N�[*0�	+j��_�/n���b.lg���pDT�pIE<B����Yz*��֋4)a��F�Al⻓��j�����)qa��BZ��<� Ca������%��\:�!��{�]������@΃��[.���	Vؤ�9uu/�
B�(�� D���W�� ��}}�m5�A��Bl��P2����<��� �S�bn�vbY=V�[d�UxJҒ�_��B���ф(�����]g����p�σ40����}�7���%�Ŝ�i��َ֒�����y�C��P����|�Q���)ϫ���h�����>T��*"X�ɴ��]��[�*���R�jsm��
��Ү�үF<ݕu�'@;wr�������a0Im���;� ��������O)�]m/W�����;]'�j�����Ƨ�	Fw�jT�)}����U�g����8�Z:ͬM s�肽ͳǳ�(��,#��T�V~;_I��׫���)��<�6ꅄ�� {�?��@\�3OE�.��o��)��Ņ���l�����a��C�D-����pl 
�A2�>�<=>�y�<ͨt��zV�>��5�e���K�ZA��z��M��AU�>�00Ӊ�,Z��	e���]>,���P4C��<_5��G�(��q�>�|O�<:����Ln�%�e�NҔWP������ܬ�pE�TNdQ�K�JX�a=�40n������4����˪��� ����(^�)2�Mr�JY:�����l���B��f#�R��n>�E�v-�G�=WMc�A$�n�����P���9���TcLC����|��)��4�[e��k�=�P2z�O����V�6�d0W'�|������?��^-�s��X
YG#}�U�s;�eF,B �6�N���NX��%�2��>٪IA��Xf�;�m�s����ɧ'SganfX��Ǎ'[v����8��Q��q����� _��K`�(.��`	��1%�\c$��n.C�0T�ш���g@C"��7>�T+8&�(�x8��]\�X~���[�Ѻњ�����J����M�F'���y!�Q�n]��=�؜j�.�]���U2	��s�T���<>�?�'���O�)���=�x)�Ѧo�Z���5�
Zv$a�Z�rK|�)�4�;�I�:0��9(��-Z��D��${�Y���)��J�Df�F+�����^�T�5�L�)�T�?��S��|Ɗ!'4��*�2�OwC%5��h��4���&�ateJd�5HǘZXΡ��eر��>~ܒ<�!djo_��]S}wg�T=�h�+�ե�<�m�A/��w̬�v���.�i��=E>�G��2D����B;�f�1��Ec��!�C�Շix��*1+�;�nq�Y�h+��I<��1{b�� �X�:z0H�'���f������
�]�ԓ�.̧Y��OXė���d�R<=&d<��,�A���������'�$6tnĮ��ע���,6D1pJ����''��RT�9���" 7��'fE@^ѢE�cYjtʖچ����,����H�eF�la�Q��#!\���0#��ib��*�/��:��{*�41��t� �d�F��<_;�U�̵q\0�ͳ������~�~P~,�!��Z��8y�r�Aa�|5(�@�7�#M��	�����8���71�>N��1OHbp4ue! p�N:�
�9�_�4��Z��_K�r���{�\�SF+���3�4�4��e����n���[�׃Ⱥ{�
�7u�xb3L�_u̧��R�
G�;|~e3��E='���/�\�(�h�+H����܏�
�D��P���ѼC�0������B��CD?���6��Ҫ������S���A^
/���3|߃�y$]����gr$R5awɖҐ�/ٙNv�Q�2���g��)&�t��'�д�(�2�-&=3���z~�z��6zX��L������QW4���i��/�T�q~��xD���n=�%G�(P�#&շ$�U��
</�;A8�������0�G�+���.�
˷��-���F��"���0�/E�Y��y��WN)*蚼8Dd�?l��끧�-�H�=츊���¶Z#��JV�;��� ��v������$Q�_�A�`Uӊd���|�zF�tm��X�Vԇ�$B�Gu����+m͵�C�ԥI�(V�E6m�Sԩ���Kfɐ�Vys���� ������VM.Oz�������Yyj�f�Wu��mR :����Ǻ����@&���%}�)��)~�9>��h�J��������I��P��O5 ��]~DM#h5��N��'d��%Vx�di��c|�hٵ��/���^�a�W�i��e48o�oj�6A�.<J����M� V���@@Ք�	��ޔ1����.�Y�+*�06ѥOV٣�g�]a~�M�ǝ�A�c1�s+���n� {������;�n��f�X� �𬆳�o��]��2Z�뎶�R
D}�h�9>i�o/�Y%�g(�WT�QP7��'>�]E�]���讂��z	$o��i��izJ���->�B*��qI�����f��i�Ǣ����d��ҽ��sο�YQcj�#o��vR�h����M�;GL�M޺U�/�5���FVg�]�5rnhLI`B0dѽ"����gz��T�#�a7|Ծדc��v�/}pr!�|Z⎛����i�>�_��6[���j:F����gQ503KH	 ��G�]�t����PlQ"��H �n�����b�=o����kqf�|�}��h�?�D-j��\��RR�ia���