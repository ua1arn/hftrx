��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�i8�>Wc�#�?�l��Z�F3~�Qp|��:��pIۄ�d�
��&��Ađĺ�M�����2�m��ahdH��I�*j��d٫_u�>�ȍ����"�+�"�sL�ĶX�r�
>{X�oQ;e.2�ζ<F�HV�5�D�Ms.ٶ�(�*��?��$ck�o��Dk�g|Z�Ԛ���S�3���Htǚ��;a 9������;�1�� �a^��6T�����?U�`��(�
c��$4a���IR����V��{6�sDA����T�� ��C�T(�[�L/�������o1i�?[.�	�Y�1�q잰�S+��ȟh��d����'��TR���g�m�A��q����J�Z:ϼR:;�R9���ŉ�=������H�����y9��n9l[�U�T�6{Pd�K*����{���Im..sb�(������ԯ͙��c�/t���a����[)<�3�
�c�|_��0���g�VPj�*. ������ro� �#��&T���){�u�Vq���}���9k������DgA�]x-���x;;wjݼ�ZQ��qM��Y�Ӯ��~`y���D��u�Âµ�`Nڣ,�5����H&��L{���l��q�=ԉ�J�䔃�ԌB3q��=;��sI��u%-��������Yۃ�x����g���'�tm��W��^ҿE��E�t�H=�Uh��4B��CDХ���5/���0-��~n���F�����ˇT)Ŋ�����VAj��Q4�:�ʋ�÷�z�Wx~_<&TW ��Q�� �y��Q5G-�1=�0�'ߐ�8��9��@f�U`{)��7�!����hy��K/NM�\�o�Znw3B|/���*T�ԡ4d�DC�[
�@{��~WNa��a�݃���~=�K�p_ >�H"�S�e��%��?�noӳ��5��x�ߢA��|FS{�\7�G�D{��&���f��:��@*� 3��\Ս�\ĕ=ȇX$W>�Q`�:�.���B��|n��0:�?gP.�YG�N�Ȼ�_ή?�:f+����]�>�L�dzԓidk� {[2����Oq��cK��RR�>���uB$�B��t>A�1L
t�[��nΰ�G��_|T+jLuA�m��{�&�XK�u@'�8��Fʂ]��Q�;s��T��ל�^o�B�>����D4��ԓG�6��_�#-Q�Q(MF0qx�觷^�\_|] �� ���B���ĸ���c�`^\�2���8������V��bD�3v�c�T`,���	 7$�43�,�D�~�.�mF^�`);��:fH�a⚅�cS�>�Kq������dR����X�("c\i<o"0d�3|��P,cY-� �6������]<��Hj�T��h�3�#�:x�V0����%�E��13�z���ɟz|I�g�O�2��������S�b�Ֆ��o��ݴ?q��X��bH,�H�G�Ǐ���a}a�0ԥ�H�O���gOc*���b����{��#b�4��;�[Ԍ>�Ou� �t/��?��qC@[�����1��}���%��v,9Q�B�"��fT9*Ί�^F!yx�w��7�L��z;� ���I���
.�4+X�4:Vx�����JL[�ݐ�ߥ`�椳J��	���$�Dq�|]Bԓ�R
�/��L=���%�8�'R�fE�r��_v�(����p�l �4J��ȁ��ѸW(��3��"��^�JI�q4�����O�y��%v�q����6�����cT|h�����aZ��F"^>%�o�=�g6:�k_1��7�|Ҩ��+��9GI�תP����.����4���S�Ѧ;��֖J�ᾃ�	�j�;�``�Uw��0�J ��(��8])�Obu����R�×݋e'��R�6�H�5�G�D���T��
��[�{Ra���T��e�
*�����Yp��{��(_�_[�R�������%���m�{�o�'�4�
�`>�PZS߈�"XH��G��z΋���c<VeCγ�G�����z\��6���8l8>�� �^TrCe�HN��1N���p��qv�7LCEE4c�r��Pri���;�H��`��4����cWK���f(�5���������D�[����	�9�U�W���F�3Ȑ[f\\ϑ��x�-J�T�59��x�Nl}Q�����S��-/(iϽN���,@��������L��eѲ;x��w�Q�a��kK�ˮ[��",ԥYlZ�r�i���P3�-a�`20c���e����#�H��'�z��@�h���0Y}�wV- ;�K������S5uIa���\��R�|���6�o���/s�Z�@�K����k����ޫ�����,�?����q-u��`�ΐo�>*X��>���}��k��Ey=0�%?�2v�G�A3���fAiP�#����U�iuh�<-2���'�e��������o��ɍ�tO��d��
���$�p�Dg.kY�Nzt�I��s�%`�)�H��]�ʄ�?p��D��I�F��c0m���,��$(!��ju�sA����A�Z\4�����C��v͂a1姉(����+w@	��}*}�S��I�A�w�,�F�G�yG ��.`�.�)�ׄr�Z�M���6sC���C;_|�@I`�41zSgz�� #���k��EJ�,.���y��}VӔ�Si��m5�R�O�ʆ��ZE��q���FK�PA���I�9n.��o��gT_��$�V!T�0��|nkH׏!��آ�FR@�8���"ƥ���%,]0@�6S�G��2Z��F�VՃ��6͡HF~�C%Մ�a,#�1���L��O��7c8VW�{b�"ǒ&��蟀�Lۆ�Y9�� ���7��Ɩb�JJ��X�� md����uT�ߍ�,Ѩƕ��"y�ʅ���+��n�e(:�`�15�F�݈NBw#������-�rh�C%�7��94�� ��
��n��|vҌ?�8�_�/�)��KY�l��̠I�=+�卬d��*��0̔⢜b�E���ֶK%E�m+f�(v��S�x��Ɍ�=b�2� �R��B� C�i�HR:0�L!"�2��� ���2�%��4`8���U9w��p��`��凤�����B��'���W���R/�y���L�
��JșBv�����cړ��!�T��lA�@Y�E��yV���hxY������4!�����s���-�{_��h7�~�XK)�xYR���}���R���?3p*]a������k�z�K�D:��U�=�������i�b"Z������x}$�D�g�\�w7ڛj//OEj6&��s���ϯ��y�{*��|��������]���<��?S	���$\L�}'�v�I	c������m��够�,#Wp^T�Cy�K��U�M������>�x]��[�}�(����|ZZ �:�
ST���(��j.�F�+��#�~G^�����6�W�/Դ]��J�"�U�p�֫�Cp�K[�l��G��k�٭Q����, ��^v�K3�'����i�rg���"�!'~��)��O�[bI�v�0a� }2��V>��k�Fn�:P
���!���:�����$k`�x�T8AkX	q��H��H�=��;ö������"�����"���.���m �k�Xً����ƌ��p�+P�͡7nZ���,��( �af#���B�� �r0��<��?_y8�$�ۆ�ݞ����,�k��e_�"�BN�+�)y��ٟ�G Y,H�:��(�!���@�=޻�-d�bu���eK��1g8��Fehc1��R�짹heU#��Zw�`�^X��r�����&Ie����v�0����\*�X��������"ZZ5,k��#��Wss7�7���5�YE�����#�!AЫ�����0mF| �ѯ�j�r�gQ���	f�	!b�u�lNZ��b���7	��tb�M��Π#l�!���8�q��9�k���,�V_9G��e#R�P�8�y�E���ۖ�s�vcԵ�f4#T��%X��խ�Y_g1\��g0%}cK6{� վC�Iik�~e�2�L��#|�޾9��˖Y?AO7�:��#���c������[�٦��9��`�iI�xd,:^cV�d��o�6��k��#�i�m� ���d^����T�L�كx��(R���C �Y~�
���el�Iq�<|�Ғ�c�J�|��A��uބ���_W�f���JDBΘ]V���eQ�c�@p'6���z��]�n�L���|��
�KN�Kq�ds:Ԡ��i������Ƃd)L��s��?zI'#;쎁"���i&�><����{�@w9u;)0��Y#�V�Rj3ɐ�l(��e�z�ӭ�s���S��V�-X1�i!�g��zZrrv��>/$K�(�S�h���J�4k.�B�-�
瓃>y2�v&ǜ��&��1=��S�{�V^�,���,A_�}����r���EI�v��[�/}/rX�V҈�(�Ͽ�1�tu�
 ���,Χ��a
��V2u���7�Êί�Ga���>�1t��ͻ��0��RAi\�8��+��dW�5�҉տAeoP����	�0u_ɴ�~�خ����M2���|<Ѕ�*0#����}X}�=�P��:��G�;L�QB:���yt��./�g:[^C).U[2�>.sJ��߁0�7oS' B��kТ�g����#+~�c=胹\zC���������U�ܧ�%H�Vg�� ��$Mv=?�O�IV�;�-�8���h@�@�7	k���t�'�L�o��Q�y*���_oܵ�x�sW�!�6W�X�N%RFq;���к'���0HW��rf{�~;�4�ʎ3w���5�lT�T�L����^"�h�q�3�����Փ܊e��P�s�.�tMj b�9O��Nsd�����R�&�2'��IŊm�G�����ŕ����N��K����ӶG�'O}�f洈�������`�\�NB�xj��Y��V�_H=�g����c�'_�Lf]3��	t���!n�&�3S�1�g�m|���T�x���W�kg$3;t]s�j�ƽG�:�K���ES�n���.�eѯ�ߵ����5$�偺T�Pc;�J�m��6�Z���?�V�$�o,��qEg���z��`
�J��u6
S�5f,S)�B�m��eI|E1L��Ho,��ٓ>Q߃yo� ���d��V��O���� �#���T(|n��"b$�pW�d�8��I5�8r��q�W�))ުԼ6�g����}6c����ba�8�F`�g��&8)�X�� _�A)2�2�eL���29�Ď�7�
c�;��}Z&~�U񎁣��d�-^�y">�%�.!~�h=�= �T����b��g����Y����0#��A�ϛ}F~$A��va.~�����P�l�E~9"$�*�8�g�̙*i����
^�o6tii7:띱��s��)�)D�����d ��LQLW�D�.x��`���f�_/��[o�΢�L���?D�Plm	�pFը�O��XO����s��i;� \��!�P�������^�(�Yjہ�9?�3
�l��{�S����S