��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���Y�՝����@N�6�-*�2�wb�-jv^���oeT.C�j(~j=��	I�ҵ�Ӟwz���b��c�M\o�e'�l�� ���>L���}P�Z8kն-\��"~e�$:������ ����_������2�2�g9�Wc���zF�!y%�Z<��Â12X|k��������4-��w*l�Z�fJ�#���N�V���,?���D����� ��	N�z�LӚ����	�����?v ��R/�O�5X�<N���B�6�X|~8Km����T0�T��*�2�᧭e�J�� ��2�K���b}YW+P��\��d۞9Nl?>�� B��Ut���h���(Z'uYC��< Xt�Qb�O�I=Ń�U�o!;�O�a9�����v�і_��u�䐁βZ�zU��r�<e�U�+X\�VՈW�-���-�p����YW�
oN�K���2Bw
���}l�{ݟ7�A��n��L�e�I��E��:\,����Gu�y�a �N5�Q���G���/�{s1>��	�^�c �ot�_]���br[�����������W��Qd�O��[������&]~�N��T~�fh�W�!a=;`i��r����bd[�w����lmy���:�+�ԔWg}�T�27�!r&+��ιVwB=3�Pd�c ݊���f���5E,z���j~�ua��^��D՝�g��r a#,�oa&�/�Y=1�8��Uj�DhçZ�i���]�tO)�^�.�l�  �����gO��,��ĉ�����~���]�{D�O�!�	ྫ�m�7�7�k�⍶���5j����&���-�_Xf�Vd�!����Jc�?���<�zi��x{��;ʢ-�+���-�@N����µ�N2���Д��k��K2��E�tu�y��GE�3����Ɗ�v��������-����j!#�ˉ����H��f݈���L��-�5�2v�;G1��l/�G�}pbN |���=��ѩ#u��I��4�|��}���w�t'���pm��R��c��2ʅ�q79tA�:P"��3�;\�Q�2t{�&��Q���a� �:Gb_���hߔ��ʓ��yL��k�*YٸUS��3"X�!Q^�%�8卼i�Rw��'�;����"[%���7t��j�^5�OP�G����3�+[���T�"����c��5��o*k����y��ዚ���a��d��!x��F�u�V��G�-znQF8��;.^���6��x+�j<�
�H_�����\d�����UvSB;`�1T�\L:�h��)�	U�.��#\eҵ>�쎔�,YǍ���p�F�H�iʑ�C�e3�?Wx��|_��j�Ԩ�d`J�U��sEs�e���������E�ƛ�ɟs�ݖ��"���W��y,��wu����sup���n��
��6�����jQ��>K3�j�>�L�' #oXF��o	C���F�/#ϩ�	��)R�E����H�i�����W�擫���;R��-[�4��(�w���,��^�MBKBYo�u����S���u�ڽ�d?&sG!/��ߌ���s6��=/���hL���Ǖ�c.�G`!����P��\�!0��&��� ����j^���[����J�m�����r}�k]Jv3b�c��)�BI�t��Y������K�e�+e- �h��x�=Wз
�����+����[,��0�:�`��♨ʗ�9��b�AgQ!�T�؋�lw:�
հ��%h�F6��a���E;�w���O�$�!�(hd���w���0J"s�dXa&$O��siM�eAY6�V5�WNL��=��s��BxZR�(����FWb��y�����t����M��Mbd���Q��J���O��ޞ��������2D��L�{�`j�v��Z�lK��HyF	��!���W�_�!PE���{}Dkb���5���lD�Y4y9��Q��v�"}�X�>�ʘ�ZE��1X��==J|�D�o��@ɏIa2*z�ˤ�n��>��n�
L
n��a���#��5>��3Qƞ����D��	p}k' z