��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b�8N�b��Q��|^6 ��Ӊ�}���.J�Y����c��W`E΍2/v�KѨo>�$������h�f^��/�-��Y�F����dV鉜��z�w��Ę�H�j[�0�n@���07��?'�ҭ���J���l�@r�b_{-����:P}�]:	 &��5�{Fu9w�K���y׉��Q�UE^:@o˷��!?h��}��IO��М���W�r�jH2�k6E�"�AG��6��8L�M-b�Ǉ@�6&���]�<9�竻�n��uT�t]�(	˝�y��6�2䦎G',!��mK�<���n)�m��8�T���G&�[�+��r�_���a�J?zHvr�qm�V�?�e2��")ϻ�m���Ch5�.�p�%Sz��TpɘQ_ס�,/t�Wm��y��!3�WpJl�oo��PDd�׈�ޭ�Ư�Ζ�3���k"5�ߧ�=�
��!%����6��� b0�Sz�|���	 )�L�~��4*�`A9�Jc�k�a=����O��v�H���h���=�S;:vD����5U6%���h�}�%�����\���ӗj����k���;�g71!�b�*奶\ٷG ׯ`���yK�� �.a��<�~�괤 ������F��1th�pӗbi�����Vs[���wK�
�c+��Ω�1�����]��#i��Z	��5���0��,n����/=?9������R9�kJ�ѝO�c�DԐv�	�[�uvcV�y��	+�ˑ�A������wx>m�;�9Q��3�^�j�W^B/,^KbD(������Ŋ�/g)�{[����T��G�8M�t!ս��V���hm$�hI�H��6>��+6-2Q�=w��l����7��JW�<�{��R�]�/,��pZ�'4@V��S���>7ʯu�ˆ4�!��ˇ@� ���n�rp�N�p�	s?U�%��5S��߼��:�@5��?y�L��e;�i�+��l���	/�4YEt:Bq�-[7��@�.�M��_a��UI�m7��ra��|^
P�T�N�j}!���KɃ�e�����[�N�A\r���_<���_;�j E�y}�C͖�3g��&	~@��[���cq��7�f�Ƀx���ޚ;�G��ƣ+�QŌ#��u�k|-Ǥ�!�kP��e�uY�۳S/�qГ��o٪�v���Eͦ� o~���k��-^���m�ˌ��Z7I��WuVt�S{K��, ��[��?ӀٸV<^�=�i\�iwZC���p}9��C��3Uq��ET�.�U�F엒͸�x�[	��*+H��Ld��}d��Tو�"P�Q��!���e��>)��BJ�8Ӽ͝2�Ǫ<v�B��P��p���%"H�;���XY�P�佱BR!�&���עq�������t��e}S,�Gk���D�q��1��3�� �|�����yo/���IiUB��.� x;��� ����Kif�vA�{�a��m?J�l��當�(�J�I:#s�e/o2������_/�<�����U�C$�݈V���4�V�%���\,��X�w6"K�
wO�3bJS߷�-P����W�a@K--�nM07��v���>�v�aÞq���'ߐڛae��æ�0B�O���d��H
q �(4��X�� Բ����H�4zC~Y0��Fq�.�W��i��{R݉��+ⱊ��O�6zn�6�C����_j3#�G�WlBp��gϪ!��C�ԯ	�JWG\�J���G� ~��e�@��#ۖ/H� ��:N��(p�_5�?��i��.�k�bN�����}3�\�Hc+��vo���Ն�!_Mm|��ഫ���`��������F�[o�G\��΅��S׬��H���1�A.H���h\U�>���%X�3D>��
=@qc��_��ȧ�c�0��d�4<��%�a^���D�5��{���]��n�����>/S���F`�B-�m���3H��Hv�0�W�!N0��e�B�����"��5����e^�\4�$Jr`}���� #�!�7N����1���5�����c����ST�i��J�������q��c��H��Mﾦ�eJS��7c餳�������!{�i;X��7F��R���Ʈ�)��S��`Cz���ط��C0�`3@�Ƒ�=�S8p"0(C��k89��-*��0�~�B�B4�����ѷ�DRQ��`o=��`�Ig?"��W��~jgs�#�����~ak_�j�Y���3G}dUD�|�3z��<S��z�wp� Sd����ϐkm��g�,��0-�v�\ے����|up���[�r=5����Q�$;��\��T�Z2��R���~Z���6�;�HX.��Ugm *Fr8vݗ�IE��t�Ny�v��$rr�� ���9^%\i�!�ro��0�A���"J�
��w9��,����t�e��O�d)��US�kOmX��4L�}�
&�k��٤�˥���d�l�Є^C�6��籒_}̰�qH��ul�V>�3N�'.���D��Sg `mf���[�b�9�!x
 Π�����hV�����V����U���~�npe���SǬ������z���1݃Q�t=j�/qu�bq�ag��b���C��<���krE�����
���#�[pP���H�ԳR�1IP�����i�3fϒ#o܈��"�f���T���C�pcҠ��*H��^S�\ GI?ܦvf��/�zp�zZӭ��;<����9�c��C�NW��T��(s9��/��7� �c7�8�ZE����o�~��.s�����2_�����+6�ĵ7��HDd� �P�/;/o-����)���V5:���i�U_�Kd���_!4<c�h��nj���50�ܮ�l��b{�M`TT�~���p�����*� ����z���k�X�؊�5�2��U�U��E`�D��P�;��sǉF@��k�@k[L�coڗ��� �m�[����]�:	�X��<=�n\R�K~����,S5��2Ԯ7�}zS��|�4���˝T6�;aZ�:��S7���\xgV����t��\�l~˞�c��oP�:�RZ�@���;����z��Gl�YfFbF�I��\1���b��#���3��}�=V��rC�F���X�!'�-���>��4���8�Ҍ}�ؗ�%�/dADk�<��Gs�r�Ѵ����z=�֞"��X�P�ڹ����%PZ���~�#��?g�[�c��<�иF�ӳ�~������<n&{�J\���$��KGD'��V� �a���ۉ��N�O�S �������/t�t�qϻ�ȶ���
eQ3�R�0��փ�u�m?_%���H�Z>p��I_����}�|��m����*օ��%�Z� 5d��#��!��`���~H�닗�y��鄺�Ki�����H���+S��B��t"�lS3�;&�9��̨#e�"	��gL��5���1����F5�,r���د����'6�&'��x����38����T��s�'��<;������c=�pMt�����؊��+�:���r
IZ�"�ܜ(�ܚh�)���bY��r1S�x��ى����.�����PU��M�?"��Q.n�L�{�~x��<0�0��o�e��BS�چ��~��h;T��"����FYB�!i�'#� y�jz_� 3՘�'Cj�.ep[�İ�ߏu[���r��H$��$�����=kbW ��Y�q�X��"��gT�/���G�E�_��뽿�Fj\�o��1�sM�9|[u�G1���M[Ӿ�sʝ$���ٜ���@7��l!
@#�m�>�� ���G<����a���QR��:H×薢����a-=��%�RZ��.���q�.�m�UY8��p��&N�B��&'�5� ��`�d#�J1T��ܝ�]����!�gm,��>�����F{�?u�R�>�����
�'Gw���A��)����Ỡo��^
���=	�SI���U��ۣ��M&-5�A�����<��8�-������f#�3��ܧ�2X*a@+��ؓǨ���)���p_O����	�뼫�T�4�-]�_|�������,�2����t���&�����k�1 u#rI_�<��6nG�+��(���=D��������Z ���N
�Z?�8F� ���q�1
Q�������f��2`�����[3�	zb�jK�S�H���WLw��c�T�BO��X�I �Y#��W�&��[�wACY�a}�-��B�|�.�5R�̚O��[��Y�2*ΰ!B���`ZB�یW�:�(u�P�xa#�W:n�x-�Ս�D۝��r�ϔ, /�။.�p�!k�"�x\�����I�LY���d>��9#�i��+ѮL��,
ʪQE���iY�>���ߒuܢ���_U\��]0(��0l�.�[ԇk<@��*���O�%\t�%Mw��ܗө�'W!=H���Fz�'c<�<�ڃ�lu��Q�����zhWD��l���_�����i08?�6�)��Y/�vtd�9��^*���3�[T�ɨk,T���2D�Kl��s�НG��c�_g��Q���H�S�1���[�r���0��*f�\���Ȯ��B��4V�o�$��x�b�)e��WJϬ��<�Vo�X�a��Q:V�� ��/a��8�����q�j U�(����m�u���NZ)nCb	��T��nbޱ��J�W�I�(�=�Sp-O�����ÃH��=OÆ"�=44���J6tF�k�o���,9����?-_j��}��˗�
I5�΋�]$��v��r��n3 ��b3N�~.eM����3Ea�Ar`��/gF�Vw�$.<���.Ģ"�6z��?ܮ5�n����c���*V{ ����y�V_�����xG��k�l���q �%;�}~��F��Js��������{~���
Lv�
G�d�5��\���I%\�s?�l��;����X<�6T}u�k��Ϫ�XţrnG�$��x�ǹ/6>�H��pl��w��(�
M�y���á��,oJ���Q?��\2�ܿ@�d���f����|e�#����k�Qͱ��B̷�0�x�pdf?��9�wG��%B>1���}�.s3:�_A����_�Dvd´O��O����B���wp��Z'u���V~^����PH��c,3YDߜ�t�!b)�2��C�kl���k L���BC@���S��ҧ�h�Ha&�Yα�N�Xt��#i�wL�[��`l� d!���v�޽���C�d,��+ە����C�E�q)A����?�F%bo����!�U��L��4�[��(l;���H"{����9c.=e�"��G�9��t�ה�m8��e��ku��u1ya"�ہ&}@�l)s7�O���,B�T�@$�کB�;Y��4� ) 4��uPE��aiC��MV���)�F�A%j�p���S���}2�Ff�A�\�M3q��	�
wm�i�wZ��|m�:=�z�`���A�Sx��)�� �S�����I�O��[A�ߜ����γ PǓ�bH���q��s�������"A� rߧ��BZ<6���F?��i��-��ֱȷW���xy�_T�~\�0�\�4S��!�ئͅ�U���Q�s�m���
�87
`T��*���_k���x5��OwD����g#vp�����~�j��o�O�&1ƽ�\1�6>]�����;1��Ç�R㑽3��0+-����|�)���J�3cs�����BjlrY���Ko��N�T(�fb��`��N����)���B��\����A�/.��-��i�m+=s'�c�������~�C���|�c^?����VQm�Ư�r?X$y�@�,.	Q��P�V�fE����J��n���b,����شQͳ����#�F2pn��D���5Ǜͫ�G����{�"-��x	����|�	�� y�#�z4wjM�nj�r���	�h8�S$N'{�'>b-m���2<r~��:�����M	$r�>T;#��]�
�
���[a���h�tz	$Ў���r�$�E��� @�3��٪w���f{��R�����ȩ ��Y�Vy?�q.T����\��zB3�B?�F�YlNMϱ�(���+��LU�z��ˢ%|���
h��H�OH�r�X��]�1ݧ�����$��T}�4*�9d%^_I|�O�T��\gYܴ��T��tۈ�] �`�D������#1~��N4�>�sB?�[��|��!^��(%�'���I�+$`L�*��/d�!]�G?�wvN|�$�<��u �����-�Ꝯ��g-� ��3&� ��:���O��?%��������� ��C������������RJ�B�����7���.�<�|��w'y�[S;C�L���ٝiD��i*��:)_���F�e�g�hfcj|N���ԫ7=�g(2@@3t{��i.ɕ&�����*�
p�뢔5��
�o�����kzB��l/��.NC�j�nZ�^�w�2�i?ۛP�c�CC��g��/��YY�C1���.k����
<%x0�Pm�O���4����z\p@�N�m�r�L��F�|'��?�vUȝI���ԍ|;���ҰМ��y� C}ñ1���� ��S���Y����U�U`���Gki6e6^^2�9a�I�.���@��2�ĩ���\�'����������$wBUQȿ�&���m��vD��J7K� ����t�d����&+�l����T������vmC�G-�����!���B3�Cmn���K=>��m1T�,Q�γH��Yn������/���N�oA�ܽ��mleGz������ݬ�j�ti\BWC��u�r���lp��w$�tHt�@��(-gt��`}��gBS�9C�D� T@�*�U|o�mX�}� �L�� 2�2�5�~��"([�������~D��"c$�K؁�.7W>gTo�f�v�uf�͹����V�ߘ����Lu�sa����ҍ��p{��k���bq*�H�^���J*4��8y� �n𮌖�|'n¤l��xL���gLD�����:�X��ɍu�'Lg�X[��U�Uh�2�̆���J
2�������z�L���&_�H���#�t9��R���Aa�I��y؎��f�4�'l����D��D�&¸URmsnW����A�b�ѯk�ӊV<
�2	ݴ���6���ڦ gb���c��U֏d{����uzjoW��e>iT�CK�r]��#�[�Ѩ����L�����LW��9nx��P�������BT2������<�]�L�����./����h�e���t�u���� �5��D������ٚ���>�TPW�JXY���O�"o".M�0�� ���]!�é�*;�a�4s@#{��\N�!.����VI����0~)}ω�[��~��� ���}�{ɕh�r6�UC��Y�z���ޝ�(_�ꕙT�4�l&j������,���ݞK|�D�<�J�*D'�S�!��M���bGSK���iJKMP��7y���/> }�EZT�<i)je�	��DhVġ��^GQ?�b��W:VF+��)ӯ��Dj�8�[n;�ڐp�X����~��u��p�V�FO��&�=N�$�{��ُo��!::	E�	�*I��f 0;�9P�����+�O[Ru'�����-��F�+Y���z��}'��1�3¾���+'1��	�#�+��q��w_n�KP�xJl���@��Z�}P�w�,�>T��5l�9-�}���c'�Fsƴ�(!~�=T�7��rM"@���>A�Q{�����X���7��%6W ����n�V)m�z�e�s���ַ�.4~��m��ƈ��zf�@���h�?�GS�6��e�d��u���1�&2P��^)`�ӈ�)쁦s�*�.�(�F+�;����{*��,e�W��Jl�B����qV	7]�>�� v��zh<{Cp fP�C�]9�g�"�+`$�t�|�p�D�s���%�'��@O�U�&;(��t�=H6����?Y���#��T����y��'�g��OJl�����:i� �9 }%�_�o�!������Wu8t�N;�-�J������*�&)�-�q0���R	�me���r��O�������"��2�NujC�p�s��wˠ<��*����Ga>Ϣ�,sC*�p36�~ �����?�s�k�t��+_(j���IHq�ᆤ�<dƯ+8���MΏ�j[���%��A��Ƈ������W2|DЖ)sY��S��I�1����� I�6��[A~�y���#�輔yW	�U�����=1��E�=�ld�w����C�8�֔�E�5�PU�Mq�X���VK)�aS��O���B���b{^ֹ��R�����ݲy�f�x�Kk��G| ��p��{�n�_�֟�� &��R�4T�"���r� �ʔT�͜D�b>L��a�?����Nl�o�!��VQ���l���v�SU��\;���~�
���q��Z�D���S]��1E:[c�+�!�c��	���9��;��Ҳ��������v�(a������Zuu�D�5���g~%w��o��Q�r!�].6aP���m�����˘���؃E=��!{��[�1��T8���&�ҲQ��M���Y�S�]�%%fU�fs��Z+�s�8��ov#�Ϩ���{��6[(�̈́��z=�V�쐢�f���ϔ��ҋޡ��c���;��ٲ62?�0o��4|/�U������U��aΗVa�.^�_Ɍ�ژZ#	�g�3	42�D�n&H&������>���1�����y�L?��>5�fo�3�>�M���5���N��`K\�%�1��z�R����k!�嶝��ހ3jW���ƌ\�a�����H�����t��v����tj��9�����Y��h�� $ ��\8t�0y�ϑ��~�$w�7�tT!UF"bOAj����e����s��U͒jP
L���zh	)�>�������K�MvB�l�-�?�8����Qف� /`X�k*H�R�8r��at�9�����m���;�CWK`1�D�ڽ)Z����o�W__c�w�[:b����mBz�"sFFܽ�_��~[���RH���~�hs933�2s���A���M-�%��Iq�F��"	�;ɵ���fc'@p�����y6[@�6V@C�em̴9���ؘ��
8Tsg]z����y�=X��{x�� �E��Ye�B�vU��5�M��Q ��V@�z�����T���F$=;�r�>{F��"���p�n���{m�f`��H��S%�p���[��&�5q��X0�Q �+��f�A��t,���k����"aw|#�������Su�,�ѻ|!�2x�,�� �'.��h�j�q�X���h+g��q�7��vj���!�v�$�f�В�V�w�X��C�/�U�0��b�`����K�"�i:#��R���"F�}�ݗ)�I��#����@)���B~�Lۜ�xAi�Ð��7l��H+�H��5�R��{�/���ѭ䋇]&���'���H&���IVXr��܃�͟F��ٖ�l��y��8��s 7���9��6�4�?�Y�`D&�]�^�(M5��T䟝ƻ���i^oPz_>�Z9�$�m)n{�9�_5I�r��wL���X�7BИ���֕}G\.C��+y�R����A��.K�m�R����"�T��h��f8��������t1�@2��awA�6�(R;Z��k���f�=ϕ���e��;?�1��7�с�ԕ~������΋����8�� ���H裴p�Nf� ���M�a�jp�ƶ�����`'��� �F��12���A�aM�n&}!t�9��9�W�y�Q��ى0�Ų�6�1��N�[�k�p����T����F��% ���;��4n�\~D��J�O��3+I֌~�?�*���ؕ�?��D�fm?ĺ2�7NFS�b#�b
Z��R��ps��B�0o�3��AC�,g��?H��@���`���/͆���?e~y.3�&D\0��[ �̝[��g��bvN�^�������nzTY9�b%��Y7�衦�S]���:)�Cq�Pn�����8
��yΆ�#���n�EXт7��O	�k�.?$�}b��;�b�[�H�##���RtN��n]�H]�@��<;3هA�@��t[3# ����łV_�j`5����d���?�@��s�2��V�
�2fyɴ��|?�u݃�ݒ�2�K���fT %�x�u�J���!-��ݮ7ӯ
9�-Y�W�ba��Y!?�j�l��}r�9���{+�)� U+ţ�Ds3�碮�`�g�	��K�b+�̄։&�(o��b5��yZ��GQ_����7�qabZr��@/�y�5�����YZi��8)戀�@\�
��=��'=�UygN�fXo�(�F���G,����r��S⾮�����D
P�z@y�=��b��{�D�mv'ڋ��v�l(�On�}vmb"CoޣQ��錖B	����
�@���Sg�P�٦�(L#Ʉ(�N�v���A L�ٮg_/��4��d�u;��M|��W^�(��Mh�:�b�Z�f�AX_=	ꓶi���w�*�<� S,�%�C�g|��$q���T���b�Q A�m���>
�����0TCjj�����=�����F�����_���N|F��(��|`�D>T��1���%����F_p��3�a^Z���Ye��&#Ȫ`\����r%��<X�%�(���Y~��V�YW}A wG��Z����1�����@n�wV������.����`���1k�R�С�m�nP����7���-U����Zv/|��.b�(%''Le��k�^Lwȡ��>u*�'�/��U����x�pc��#�����}\�q{�1�RՄ��6|:;YU��ɘ/�����*WI�P�|91	j����)�v+jGi
��3�"�j�������e��	�p�P`bL�B��O�������r=9��\�bwJܒl�-��Ap����Q>X `��0�Ad�`A�a����y �zדTPe':x���{�{�t�ձ���Q�'J���g�qN��B8�벬�*����S�EMDd��0�eυ�^�u;2�]�r=�m�{�l�|��Q�ێ?��{�d�&�=(��k�B��t��r � �V� ��Y� �T�}���R�]��:�1<���E�׎���/(�I���8�(V�j���2����I,�u�; �LVLϚ��\���W�f΢�2�� $�Oe����޵}]��(<�������7迄�usY(�M&Iߺ���2���.�������+�;��GS�ӑ�n�q�|zOʦ���s��C��Yh�������47b�KB��~b��1�
`3��X�@i[>~nݑM
�h7�s&j�!�@i�uG��W`���!�T&��r�`�����&x��T %�A�S� d�lBE���)q�n;������Y�΂zͿ�� ?�8T�?���Ѣ����b�k�O���z��ۗ�e/;
q�eq|�vHM=�&����YY�by"݌1#�ؖ������S�S_��5esE��AQ&�����E �V&?��J�:��C]/�D�Όi1wT���9x4#�RV�CR4=��H0hVU��d��Ӯ G	l���<�u����n�
��M�I� E(^�Dt��CG��}~�ϱG�K<2&�z'"����/�۴�h�fݗQ��hF@*�*t���@ttFQpd>r)[��>�I�Z�WI.��b(?|�7g�'03�� �mɫ�Om�ى<�9�z_���!�{�?�WI}�(}���~1��@�(���Z�w�>:eF0V@]��Q�Bφ�qlQc� >�[�(�0�q^��B��R�G���o��؋~��y4A;"A�q�sPޑ��ˑ�g0�0�dhM�>��.H�׋�p��i�c��͗Q�c{n���݃q�?15>)�����������ڮ��6��O�6���>y�y�K��[Sw�� ��(S�n��~��dAކ��P�E��U���)>�b���d��ut�L���ĝ��ԃ���F���-7���r�ըCy!�v�F�3I]��o�8�2�> uVkAި��%[[# ����]
��iQK����cjo���|�㳿n���
��I�㵄"0�>ѭ~�ےy[K�0{M�\`��� 5� ��IWhTI��2��,���P&n�L���QM����d����s���q���qе�#�Nb�p��j%w?;�F�N��i6k:��3d0�Q!��G��%�+Y�O,O��,DM`�!�7a�T��������Vwbk�Ԇe�h������B9��v������P4��Z�+�m�����uA��Wcf����"�F��ӡE-CˌÅ�x�B��("�����m���<����a�)�O�?c�\�Ew�>��2����mſ�����M�ib�����2��|���ί�D`���(/�e���ь��	�m��A�R���Ч���N�� ��������(R��0{��=�����E�8gE�k�1�����XD˦'���D}sˇ|H*7��W(�$o�l4���ɹ���<2�渶
%�X~���8�Ȁ�5s��?%D*F�z�� 	�wB��>�u�܇�G�~j+���$���/�
㮻q{�fs��J�S��el>�5t}R�P=�=�4�`���A�ʵe��y�p�ӷzQ�܉�\nbd�:�Wy���B'�X�WX!z>�H��y�m�\6�ѭ�)�:*]{
F�V3E�6����rAW��ͤ)��&zk������Ĥ.�gYеA5��*Ri���T�˫Ÿ�g��a�x�,%.��=���.�`�Icd$�݉A�Q樭VQ>��;(A�KJ=�::�d�.�Z�ר��O6�8�Rި���~���0���!��UO뀉%����)m]��6�xX�)D�~O�Qn�����w��6��F��u��g���������|�ͬ� 3 'x <�_�>UhZ/��`^cVR�y����lD ��=��y��(�UP���C�r���D*S=�V����u�R	)\�}���M
`6P^��ʘ��R?�O��fO�4�*����iF3W��7ȑ�)��k�`�Ə���Ƹ��������i�)���u��p=vHX����%�Q�k���6砞le)�_CAC�M��!�3ds ��Y?�W��>��nG�YN�j,-8��ܛu�+h��q�c0�ù�zG��@iC��T���U�J����N0��D]���WI��]�H�ЪK�A��?.B�����G�J2^@Rz�Ίsn��i`Jڑ0��ۆ@I5*�2��Q5.}�͹�݋j�vJ��Q�~pyo�1
��Y�D�b�e �W����O=�St��)-2�Q��x����LH0@�K��&�9�}mhb�Z��ԅ,`E�~4�*�W,���.6,JKD
�ATm��o(�"^�X��H�����Y`)���Np��0s���)��8m�8�4ߝ-��K�yj-�=���RU��&T㏤�Χ�O�P�V^��.�lX3�d�t��B#�M�JZX��?6A�L+�G�ڼ���gm�������{G]�i�(�d
-)5�f�嶹mѯ݁u�1�c%�K3�����mp����/c���E�?�:��A��J"R��Ք?'NpT�����ND�Ә�oXh���p�XF>��!�,�T�lǵ�S�@�"&�ש��J�1A�@Y�)���	�fnw ��󤷿?:�a/��`���z������1�d;�@�+�h]3u}�_ �4pp?���W��6�A��tU��������V��>�A7��	��]�Aa�~9���3Q3�L��L��LN�;U�ɺ������uZ�FƘ���˛�9ϧ��bwάR��yirm�fe`ᕜ*��^�I�SM��c�l�cv�SO�K����È�],�� ��1�0����O����$��n�+BS�cѥ�H�m��b���[�1�G�<nycy�ڃ��+'c��c;O�Cך��x�~��a�<+i��1r�����k�Cz�� �ډGF���b3�UAyR��%�5��XsM�,OeY���59c�b�1zݔ͹��y��}w��У7=�p<����]>�dB|�η��_l�VR�T���x�1���m�?�ԨXGx�F�CЄz�¬p�)V�;o4;�������)�kc�Ѩ��� �F3�9��4�ğ��%���`]O�����G�,Q؊�m4XC��\�5��n�"$��)�\��Yǆ���ʙ,Gc�&t�U�N�?��~�՗\Ja����)W�UD~.�|���{�L��5��ʈgS)s��W�ކ�`��Y@��ŭ'�=�-�9C�U�z(��w���z����P��[�
c�:��K�n�	��C<{ �A�qy� M�=�s��� l��􏎧
:a�bD֟/B�7
���.�;���BT� �g��J�uU�R)-�C������\�Ŷ(�)�_�oY��G�ڳ���g�E��a2RC�x8�D!�$I���tv���p�2˒%�����ּ=��D8�������Qy���D�	_��Y|��d�j�	i���}�=�V�F8hn���0B���X��e�;e`��Qv�U$��N$w?c�&r܇U�^I]x�%����)I��4$�% g�6�'�n&��ϲuP����#�*���T>����7����|M��y=E�^ 6t� \(��@��+l]!�倫0PӦx����X�o^{忹��g�`�Jn@���I��:��pm�)����p����w���J���P
�冨GEy���O�c-���OP{`$�(��J`2X#�����vIrNNA3�g�ʭ��(�Q��X���$�'��;V*Ǻ�[�ZP{����Z|۽JhBԓT\�==�޹��4��{�"<OQ`�Y"q
9����eluR��l��7E)�X\-L���Ҍq=��M�XN����Ka�����Ih��Kp���T,j��[4�fMm��+vn�������
�����P&m:�л�4^^q����)0F��)�0}�e:HA����I�X��g�w�v�m 8~Dn4��d�VQ�<�mʰ�L<@�eԹw��@�+�+��E��3�h��G#�|	
��d��H4*EgM��a��8#ǖ%}�M�p��b�e�\���W�U�BT��u�&�[Cz��X��*��S�?$n��g#��U���O�%�h;�~� Q?��e'�1�H(�1jPي��7��9�4����q�q`6�u��gv����|}(D:�-�|3R�(�b�ȘW�!�&7X@Ǥ�GaΚ�&�$��Coh4MD��X7"�*�{.۬�w�wS�-�-hV�kVw���	�p�����I�"[j��7������K�_���$�i������jHInr �e`���� ���8���*h�]�o	��=�;A�q����� �+:;�2؄l�;?O8���ɧàI��_`T�"7	?1dG�{�Z���E8S�kɏF�?���ߔH�|/mk�6�k�����H��|#:<sx#�s��lXgҋ���Z�òe�T�#�����c���Ғ�O���7G���Լ
 D�Ɛ�hUQ���t�*Kj�1aq9�sI`.B�{�4����ǰR��R��k�l�њe�=ʸ�WvYqO�D�/9>o}��8�߄�Z��8.1w8�F��(�!���^��H2�����I�\�a�wv�����|H.�����P7ʫm�� ���v�0�?�e�L)8�*�x�	Gc"�^ � j9%���9ng�MSmo��zТX@Z߈s�C0�&�	C�j2`�H�t8�:��������BL����7W�u�d53�,ܛ�:zMy,B̴p�c�����m���Vۘdi�^k�I�^գ�wn�gB�h�stb�V��'U�}r����:O.~Rp�^ů+��7��8�<nbr_K����)�k�
��>�n�]��8Ώ�j�-�~q ��eY$-|x�v���ˈ��S���^�t6�t7�!ڴ�����5I�D����fߌ��h����PR~��0o�ɠ��`���1
A���=�`/H���x<x��/�5��HN�m��YE;
��Fs����ɽ>��5��8���g��F[c3��v�e��2Z'<b12��ȏ����ǭK�1�I�k�L��-��(&��CL�~�	x5��s�~VC(;�e+�W0��e3́/�>�A*(�G����m�w{�U�Tf�7B]�g��n��X�_fZ=܏��|�P�{�C��R�2���^jμZ���B�6@
�Mc2�!��(_%��SQ�Ef�ڧ�F���BLV;�'�KOh{���
I�����X�����	4!Ao�OǗ�#� $�x��l�:��K���LY�hFm���7n (DC��9Œ~�9aգ%�2����
�[��Lt�9O�#���[�¢ӱ/�I��ܩ<j(��@Ghs���a����F�F�$ڥ��;�PA� ��JO�^�� �bs��_wI�'��W��Et{�hT���7����c$	��6�䞺 T�2t:@�u=<�F�=�K]B�1�gB��-x�\`s�(-�!H���L)�N;� �&�����2V��U����g$]�$C��\����3*�ݡ�[	�����	�����D:��fϐ�5�0l����3?�Ɩ�i��0vM�f��v|b��=�#9��|z��*{K���;Ւ���X�!k?6�f����?�m�Mr�O�Rg�����oGB�K�u���}d:��#J��ɸ�]��%P��oX�O�j�6=C
�t�F1T6��o����R�*�K�8�x���/����<'s�����8��P�8W�U��Hj��k�)�km��i��plq_B#r⌯�4�i�N�-!��*��Y�!�Ss'X��ԦEQ�~��J}jei�sq����������<�/'(�\v�%��$|��O=mC���4�tB�u�﷝m��w���'��+oLs�]+yZ�B(ļ^�
��G�kw����xC�irbޟ��s��R��$��5�!�gI�����zZz]�����~�N�v5��;�ʠY j2�ԠmjO���IĀ��W�������K�ăYa�paX����4c ��������DE�5۠.F��2S��e-�-7�d����4yb N(�IXO[���g�<*�/�9s�:�����]�%�'�t��bP]�\�ӟ*���Mg���b���/�Tb؎��q}��	���*�ve }Z�;ӽab��ǟo$��v�Q������{+���7�	�����;��v��g���|�~��̢��z��uIB^6/YzY����CR��s��2g�o����Ì��Pb)���АF�H=�E<��aQ�!� GV��3g���$b04ʍ����s�]m��C�	M�^���F�k����3�51Ř�X��P�/��~�I��.btw��N2�P91�5�" u��~�+ci�
�!�����yψijF��V�ao�(n��N$��6�v5���ZI��b� �~>�� �&���0�/�$+��������' �fn#2�^ ה�-[�������+TA%��fǦ?Zlv�����$�0,C��� E�V����(�����zq�{z�҂��#)98��_�歿�ݵ7����|v\�怬�'��	�"���f;�d�����j>;�{�\Qb�A���t �p��en���8^u�����*�S�����Z�h�r�Z�;i� �ټ�x��T9���H�z���S��K�b-�ѣ�?�u~K^]X�Q�C�x����ϳ��KR8gP)\o��D*#��!������,�� +�OR�ۄo��wڰw��R�!;�N�5H����"�i;+�q�%�Ņ�I�ù�]��ᕿ!)�t-ǈz�A,��_�侒ګ�t.�&|�y�c�@<�8��h�q�j�?�	Z�dEe���O,��eq_v��fQ5�N�WC�9P�U���
aEP��������K���f2���ּc�<B����7�2i�s�?�q��rQ�J����#?���I������Z�_\�����kC����XZ��W��EaT��Z�����4�ov� 61y� �mH��n��Z��#�}�����i~�d~i�����~��d*���
zΪ�}���@�GKd������"����n9
o�g&��R�F�gb�C���[�"�9\�-�N�}Q�e=��5��� ��O�E͝P.�Tڴ���%�&\�!P�/x�	�����|12��!S^�Se/$4��uE�x��%���W��/Ք_ �P���!E��2׾��a�w&+BBT2�Ԃ1ќV����<��$���t �5����BX[�2������N��Eؖ�m�9b����+.��՚_�%�I&{�`�_s	�6ˎ����}�NLty��8K1VcNk�Ka�I@��i�TR���Fj��C��1�32���
��ui���59H���躧nN�������O�
Xbrz��G��@?�,*�c꺱�>��B�rJ����ڸq!�W��tP��"�b�R���	��)�����Z������J�+�I�%-���\�r����A/)ir�Zɨ����!� "<1��$�&�jL;�z=�a�����9���AF�}ФrH ���)Av�}un|h���#�g<1�%*8e�Q�gXf��m���=X��'��K������,G�Sշ���r.e%�q�&'�}Bՠ��&�:���t4e��bm�(5n��`�</Գ$>i��T� �p�&N��ILi�7m��Z`8��߬S^��>��-�l�f�? �g�P����㏢��+>��'��5�M@U�?-2�i���Z۠wk`B2����Ά����]���g�1c?lnC@k�0�~K(�D+r~/z��WQ� �]���`n��b�L�A�Jl��(�ݰ	�o�"��u�D&�;�c�?����HPkɽO#Q8Ʉ�|�ĳ�vӜ"��P'[�:Vr��v{4E(��ydT?G�ڳϞ��Gg�����D+N�����\�_0���ͱL�s��{>ͼ��P�%�N���Ŕ��~-̝Xh��+. 2+����k�O�-��u>\�G�A�(R�o�W�Pa����,�ZtH@2�y]F�3�8p��8Ŏ5����P��C��nE�$�SJ|s�cm�R{[�!Dƺ�F�Vp�s0�9L�#P��.��S�S)����f��]?���J�g��%s�ł'OE%��:)@'�Ah~|0D�� G�s;3+�A���{�.H(SݝYuiC*۽�vQ����80�dU�
��'��|���<Ϧ�k�^IG$�C��mo`sO?��;n�O=*[a�kd}07<�]�}���k���i_�*��hu��Wx��ѡ��L�\��,*������D¤�XwI���i;m?|b���g={T�:��0�i�i��<*L]@]�k�>��>��r	�R
F`����˥ ��bT����u8HQ��pdB7�s!�7>o�@�9� ù,#��y���!�1Z�`�
c���8�1�_B=�xs�~�_Utc(WV|��~�ڇM�T�s�.�)��.=L<�;4�/�W�O��4ހlq`��)��q�H�RD����䘵��/�m#��� �ZΎ�^����5λ�hxq\P�x�C���U�+q�+fi��G���@H���Yf�/��%ģB��Sq%}�h�_����X2�%�h���2��Z��L��Fܧ������5�؂ڭ��_��A�/S`�{,H	n�<�4-���8�VV�!���j	l��������d�d@:�Y*⃨��O�$��	���Il,inF�u����HH��Y�K?��]�uOS���RͰ11���� ��`�V�_S���!m�3�~����tN���6�K���ˮT�ǟ~��z�����'cs9�t��Kmi��@Sޥs,��JY"�3�#��\���Eϛ���r�:�*+={^公;��~��'{�
���H1 cY������n���'	 \�SiQ\h��(�LEO���єi�f��m���V;\s����X�5!PkG����\��22ަ�&nǈ�W���߭�s����5 ����ь�J��#�p����3���S�^
"|�X�Ef�)-N?�Oy\@E�X4��e���%���ۏ�X�t��r�)q����<���?<>a��.DH�2i�7�B0t�K�4�7�$6�.��9 0���E�+��fLnO)�Rg�Y��x� �-��4�QhGo�l�����@ij=���k�f@�~�*��-]\���kk&�aa�3%>F<�")Ф�&zh��n �̙�
#���K�f�l~&Q��]ȸJ�_���=Wz�aNx�x):.�z{�e�Ajq��8��M���q�뎬�L  Up"$��tI�eT�Mp'ʒ
�F��$"R�u��3�D��t�5�@i"�����L,��Qe ���ũ#h�ܗ'<�z|!\-���K�*�[���\�`�!cn(o�:a���x�1�a��40R�\�-��o�}K"��Fc*7s�w���e7�\�o�[��U�Y��t0�u.���?�lz���!\ �?�!����Q�)3��?R�=K`y�jۻK���Vj�J}&"{��ʩW��Yť��j����4b�+����(7"b����VB�Ȋ�jڄ��S��3�w�?gŉE1�o��)rh�!�J�^2p�>xY�>���单|	xЧ�V����3SE�` ����$�袃��'
��bi(��g�ڞ�Y�'@\���Zz��pt�.�w� Y���]ͯ��4B��@<���A��Li����ہ΢ٷ�X�m6�}��n�@SAC"�u��6�-|������;c)9ǻD·��{ԉ�ݪ]��o��iUn��-�e�y�ء�ԇ�9a���,d�+�b�P���qс<�.����4#Av��Rzg9�b�PG�8[���%L��|��K�;�wf�̃�b�`=�g��F�v�k���χ��̞BVpI\v�"X��(ʃ���֮�)րؽ6�ASrC���Q��t��
�$0�����]��/�A/��J�ٿ�'i�'�YʧH{o�?YZ����.�ב�h���`K}NY�xcH��(������f��,*�~R0������>�'T�_n��� c�a��r{�RQo�PS�)b��2����#�
�M�T~�'��M��;�X�k) �/�;I�f5�'�c�yڪ�6���35އ�Fw�&�G@j�P>Q�����L��ZZ:�GӍ6*�Z��qB�r5 ��Ǿ3�KWy[o�t�<o�d����@�˝P|C/>+6!~�>)�ِr"3��@��@��oFy�w���]Ygw�p��>��CB!�ǳ��F����~4(=K�j���`�3��xm<Iy���G٠M�T�Z��:�Y�V��p��<Ds[�L�?�.:���]�tt|���@��� �W�Z�&�9�Y�D�?ߒ�>wGLB��+��vO�1�W�����h��_��6��J�P�a��#�ڧχlE�$���N�[4:�7����͜������J�=��xS.@��K��&ڃd�lr������pt.b6�����
\��T@�+�5�:�k/	��1i��<e�n�{S�X3:�&���,�`4�}"�2.�$�e����$H���:DJ��@�| ���a_���ȊM����2���]Y�������>3��-�g-y��E<�N�2�T�%�v��y��z���U��?C��Ҵ�y/� @���o�y\�ZS���>�G���|��ڹt�ئ��%I�����X�����=YD`��lس$��tg�M�g�邵����1���RC�&�5B߈�w-�X�P��%v�氈��k$ئI� %����q��Vb�,��_�F� ��3?�N(���T�k>���F���^9�|cXr� 7��9��l�{"��c����!,t�e��|S=5�|^�Ǿ^˷��S� ؋�9���j`C� �'�Ŏoܼ�r��	�}&}v�f0��A�ُ�K4�%Lu�~��%���������ؾ�UR�)��9�Bc��2g�����!|�K0[�fv�F+� �����Pa�ѩk.��!�;~����-�W��*7]�)�k0�0�O*}�n�e��Bma�B{�)�t��y��	�~ʼ�x. �-�{-t�;��8-c֎�=I-d���mg2U3�]��N���)P+�S�2rP"�G�{5~�F�$�&��a�H���P�I4����l�<���g�j���Îz�� ��%��˕s�*vdD��|�L�/�A[�,�l�x��(y/�QŸ�tvh��R��*W�;KB���^�(�F����&���3q��:A���;N�oG����-|d�%Ғ" }�(a��u<B��3�eY��.�3m��òV�f]���!�bT����Ĉ�ڛ�AO�6r��RA{�B�����@ W�5N�Ǔ3O�\GO���������j�:il��a1�=����0-�W��Mf[d�P�x��9&�Z�+(Ue��������;��TdRq��(K���J��l���իG08�W�\ ��?5s�pՐ���Ɵ���]�3e�Q���֐���ꦛ��ޭ�r�P���Yz;X���+��D����o��k"���y���Y��.u��7Ʈ�B۝�1�q6��U0m�&X�-�D�f9�f�_y*��LU�y���Dz�>�UC�}�m~����)|(�#U������? �|d3/����瀅�����374�o*/�-I�����w��HRT�t]�D`VEx츾BWCgp�Yu��ʾ�1�Y��y܏n"��߶=��}mUcw'�h"��L@Up� X�}6LhŻ�3el�����cء��m���<�s�"�|�(֜Te�ܚ��ū�� s}IwC��ͺꃴ�x�x!k��J]�
��V-�VJO�Ղ= �n�7�߁9UБa��̏�q
u������*��'��Ky۸Q=���X��E���<ܹ�{��\#Z�V���	����ԛ��0�����u�c+�F���Tu��°<rt��/^���ӯ��cC?�����h���v��+X�#�����`��j*�]"P{X�����W�̸t���f��0�D<��g�k�@��a��7zʻ��
�-�-U2}�j�b�hOvt)n"�(*P�$���	C�����`^�{����Ht��y��$��^�-�+��}ו�ީc��DV���L���w����p�����S�N�mi߱{�GUExƹlٚ�� Κ�$ڧ�t��`���#h)�0����G)�(:n�O��Po��Q�d��ւ/Ƨ:2��*�y_�_z�W�~��v����� ޢ�3"���ʈ�;��s�~�ob�+?�c.��CGG�17l�o#M�)�h�ȝT���e��P&�7��m?ΐ.���gY Vy�m�j�LL��^��UF� �#��p��Yh���=sI ��\��U��I�S������n�'���h1čC3���G��U�@>/��y�Mx�`l�Z�x���V�fx� ������R� F��7=R/-gf�']G�_5c�lM����a�&�@���ü�2�������7��W�l@eS8������9o������l�"���-�p�  �k4��_�L����Y'����D��M2�oQi��gCɱ�سy�k_�c���kö�K��A��;�݄:��.���94O#�K�V��	n�4���Y@uV!'�L���6��/1O��C��������w�Sj��妭ʄ�$,�X��F8�y�}��*-Ӽ%���&�C�|Y���@`+ ˡ��V�B�S��-��K�3)�"�T|ܞAm�$��ߑL �A�W.��ؔ�@�Whn[�T���*;�D�(���f:2�bUBb�d�,=1"�d{���/VУ�۹%M��,��pr�/©���Qxt���8;J�b�`r�=O��� �I�-�GJ'Go��A�čڣ_�pO_<b�g/�-��Q�%�eG	:?�gA}��!�^h/���S�Y0 ʰ�N�8�����{��J\��֎��)��)�⨐�`6�X��7ml;m��of���܈!��I����L��Q�`�M7�%��0�4g�����UbTy9�E�������[y�jy2J�c�jؑ>�W=F:���?W�Γy����A	�f��2m�b�m�~r����1y}�ΰ�\6�����e���Q�p���r6[^���Ks1F�I%����ER�mwB��3⴬
{�cI���L�q������XQ~}���~�>�aT	S�/3����X��ˆc�O���U�5�v�m�kvȌ&�rM� 毥�D�V�޲���\ںM	:)����8V�,��j�=U�s粍��zE�4
]&�24��l9c���K�y!j�T�z
?�(�F6Q�h���c����%ւrN�vf��y(�＂��Wz2A+�T�N���EUE���#y��9��@r9�IN$z2Co0��ޒ[�j�f����:� n�SW�<�?�a�H��DR)AF�B�퇣�'�lr�A]PzQ򪙯˳�ْ>���*T����HY�ŕ��V�6~��+l$�P�-~Z���2��Լ�^`F�j�B\V���u���f�ew�wW�s�0��LQm���D�R�v�'���C�O2̕�2�(�M+們���M&ڒ�3��Y���w���>��<��fd�%C\�лyĵ��+����
��C9,1UX�����(�3;3R7�߄a�M���T%{0���]�Ts�}?�<'v:��� �搉O(�I"�\�A�3�u.CJ�o��v�3e�]�IJg���Ԍ06U���jD���kl�s�c�$�� �#�\�*�+�� �G�DR�c��|�@��������-
``����ط@��j�$�sh�Y-k"E5��������{t��0.�t���27Z$�Ŏ̋��|k*�l��豚v�Y ����Ľ��kگ�W���)���gT'�$p�P���yx�On:��N�2�2�83��:WcRܸ���T�RI��I�S�0����ϗh��06ZJ��[�
��MtR]��5�������~�Vj���!x�4�ݗ���C3�%��~.;ަv3�;�x���g���2!�ݧ/�J��Ǯ\}��	X�P�k^C~��������SN&3!�.8^?�g�A��$6�Se(��C���u�J��dp1����1��)}�v�5o�&�0\��$�Q{��H�+��^c,���|��{3�D�ÇI���;��G�S�>ӎ֐S�7���(���5e��	��ï0�M/��߉Q���y��v"D0�~��	�5���X�\���к�!��o�a�i���9��5���xb���(2k�|=.#Po������p�͕�f������z^�o�u����bХ��h�uFN8jA�p���gq�ud���-4"�'AF�5��٭b�=&;V�N$I� G2���*6J>�âl�lc�r�F���9ŷ�n�5,'>�z�Kq^PknQU���A�*1D�H܎�FR-"���kę��V���XQ�xZ-�Me��(�"EY��F|�{Q�p2�fL�J6�O�О�E��*!5��Z���S?G��R�5q�ך�a�f=FFj�����O�q���㱌�(3ҿ�.�,�u�D��8���W�@I�����/�A�06��^�@�as�_jm�g�ߢL��J�w��1+L<�>$��@��ʮi���t@@e����h�S yb��ˌM��h�IX[�_a�7��yA�C�Z#�D��ؤI�c�^�����!�7q!@I�@[�5�"��.0 =&zR�o�'��m��n��h��w��k�Ҩձ8ndF���ys�$c�k��Rh|�>�p����jC�,E({9<F-�'�f5�	c<tPN��ܩ}�=�dwȾ:@��Ìᤈ�jr�mHW~K
� ��ؔݖ���٦h�q���Sv�-��,�80�L����X�
D��:�昒��`���s�l�!KŖܠ钢��gQ�yV�\�ίu��
d���c�4|~�;�r� ��"t�R_!�(S��ݤ/Y����c<�}�L�KeZ�� U�-�nm�C��?]�Ջw-v���3���[@]<5�8voh�AP�<#e��^�w����1e��"�a������ts��s�z�R�(�u�	m8儞]c�$�#�ᐶWh�^�.��0m�qc_�b��Ys	���t��ZT*Yr�+�5=�K�����&
a�HFk���DY\P���ƴ�)ɻ�=��݇��|�9`4U��W�O�Cݫ��q�:K�X
{��k|����ʖ���K"�s����ޏK�{����b��B�����=@
�j��>�a�Y���:ڟ#�N�A��s
��Ҧ#�븼2>(�<E�	�leW9'O0XE#b�x3$��h��,�Udb��x l����(֙���� ��̝G�A8��6$ov�O��I�`�M�s�y������ ��_�A��k�Q��E�4��eg��Ghr����2�����!'3���鞽gc �*#@,B`׀!��=m\r�_�U���vԽv�3��d���7m���M�����P@YsG"[:D�#���9�~t�E3 �^^E:v��ݮ0m���D<�*by��䉜���	��������d?�4�΃PQ��1 �q��~y�r�y�uپ!�!���9�_h�P���P�p�$H.۰���_��$��?� E8���f 5�NtS�V����4��B.[��q��ǁ �Ԗ�����;�'���E�5?E��Q*��-z��vn׿5��S���p��:��&���,ە9O�j"���\*����Zn�e?�\�-��������[x~Mģ�łw^f��B��)�9��`q;IJV�e�k�	�Љ�}��`�E��&�6��9�^m��O�g�Jk���:[�����FS$I��6�xK-��2���פJ[�h6q�)�v���恑��t.�����g$����Q
��X���y���Y��c�e�f$��J�Z�"��+����X��vЙY{�G�	�|��G�E�g9 (8�4(L��فSˁխS8%��M�l���A_��ɂ=������;�w���LZ�o�%�����'LW;�-G$*)߫ʂU�Px�g	ĸ����E����W��@pE�GJSS U�~S?8�E�� 5fQEg_���m /�mH���10��A#�;J���١ԶW�2��އ��.��5�lI{n�d��i\�������e[�̼���eެ���˫�����N��4f��Y�!�έՈR 9�Ȱ��t�;�q�^2�q��ɜc�C�����6vM�Ɯ^X)���ʠ�S�?�����i�Ie��	��&�ř�RvT�򘰋�zX @-��1Q��I�~�q̍��?��*!Z��L�o��������(��q����Je�ʫW�,��{מ������4��| tA]��W��E�#"�P2W�)_xk���;���Dɜ�p̭2.9톎��8�����T[�z�wmT��*t�������kKZ�?�)�<���r+���G�d4={b���-P@)����q���f�ݩ�Љ��,VY\��i��� �C�9+��G����<-�>��$K�c��f*�i��Dz#�jV�(=5 ���8�@��?_>A �O9�V�x1q|p�,ɠ�Z�	���d��X7P�%�����Ta�J���3-����$�ON�c�<����b��(ID)} )�~�F�#���ׁ|���H#��)�����ilg8$賳�62\295�Ŷ�'�kC�Y@B�C�٧��j �yC��iI�Bb���z?ZQ��F�廓w^Կ�o�wD"��,�5:^ńn���!���C�(.O�%D\����+�y�<H��ɍ�LBI˺��	�5:*rW,��HÔk0�i��C�45�`ƈE6c�+Z��S"��L'���nwMQ��#�����H@�U�ޭ���:�@��)�c�$L��0C 䪌@@]���S&V�t��?%�	.V��$N��T����@�"B``6�/��ܵ���ImSL^�e�!Kh�:��#AC�
 �tXHph1�i�����D�ɾ� 7�n֠-�f�~Jj����;�pN�+��_'����mS�\�K���Xt�v"'L���?�Y��I��6�cSp��ʺ�.�z�O�eG)�xq׷��O~򙪤�߬����������}�����p����n� �hN��!Wa��7�;�@&ϣKַ2��{�"$g�VԷ�� l�ė��Bd��XA����k&��W�]@�_RUc�+Q�O@=��$Ԕ��BӐ�1�=�6SB�9@��qޯ�U<�)m��f�f�0�}���F`����{"�S۩�b|շ�m���u��F�����E�(�	2"����I�n�+�d���^�V,LB�Y������T�տ}�A���&�h���s��=�i�eUs���Ѓ���(���b�P�WH4+�u���Q�`�HG�h�Thv�|������#���tD��9VT78b�)LBe��կ�ĕ�c��_~Ӣ�1u�4�t?�a���Jˑ�����3#gL����p( �qܿL6�V">׾I4F�?��@@C���Y�|v�8�����Sƶ�F�;��Z	��q���I�p�N$1�
+ET� ����}�?ƽ/�$¨�s�.��ْ�k~���x��\Cu �r��W�H��S���)��l��N��䲩Ξ�:jǓ���|h��{_1�(_A��j]*����lS��Ω�5�'?�M�a��*_g)V	�~�ԁ�v��y�!�+�xǴ��J����qBJ�Ќ��uЛ8M�Eb��LY��}u'*��S}H��� a�V���0Ţ>��`�����%0)��<ŗ�nB���|K��@9���n����0r�kpc�ᔷ��n�g0�_LV[����B�/\�u�!�����`�'$�[0��qu���2����z1?�B)T���W�O�'@���/ub�7��ɢ�鵨�R�$��ۑ��%#�q"���k�ķ��s�*��^j�[�ip^v�l��<�Ϝ�M8���ٽoF��ņ��c�f��I��N������(�SD��tPN7��'�����
�/,,-�(��s�����6��)�\y �~�� sq��#���BkA���t���V¦e�pp�V�b�'�*49Ԅ-BCl��.rȑ�'�2�����+v��O�b����)Cj�Q~�@�����>��	��$�BH�+�J����5���D�:�� ���M��W2{�i
%5�'���v�έy���N�
�a^y\IՂ+��s���0w�'����;�D9i�o70;M谊q��]4�L�~�荫yOS\�\GO���K��0��x��*f7Ha}��8
� ��2�����7��km�]�~h��C"Ca���	М$W��棃B&Ѫ1�gdY�{f�h�wj�3NC���_��hMg�N�)wS/��9
zТ�t�u=����	̀����A]�����z:l`r0�������TEXw�6XD����cP�C�8R���e�{\�6�BԢ}��Al�$ù�}�?�����瞭d�8h�0�!ɴN�4U#V-�e:]�����ݽ@�
#���`<��"o�
���Y{<j��'���6�`��n]�~p�i��4>�6x>-<��~e���zm���*�ѓ!�{WG���o�g��l�c%1�|��>�����p���	=�*���Q��
U0��\�>7a���[l9�+6�Y�W�T'��6� �q�/���1���"��ױ5���c͆i-a�1�G`Jp���w�a�W�6��0+�}��02B*^ʽY?��*��I�u�X��I�.��ʋ�!ئ��Ŷ�x��]^40��VKA�:�3���y��i�F�I[��;�&d�^;N�s`���Tw�X	�xTk�ȩ�4�,�Y��(+�'�q�86����vFI���r�ր�~�^vw��(�1"�*%��":'�QĖ��
�M�_qy�����+����dlݥ�%$��,��Ȧ?��� �� 5A�s�7,C����҈06`�l��W'�_η� ��H�>'��1-���#P�k�	��oU���Cx�u�q��̵���$���Y1�a�1�~S�j��ճd1I�Ĉm��ov�v�Ȇ�����_ӑ��x��Gƨs��#A���7�WyGb�&�G�6v�Sd\���J��]/��\T�YJU���&���L��?����֡_��8L �D ���~�G��1���V�:��W���(�+���8�:�$�o��B�{�.���G,q���nS�H�Dnz���ۀ{q���ZY��{k)��E�X}�y���Μ5z�W��iC�������,��/�q���̣���/����e,��N@�ߑ��-�8Ϳ+|{$V"�a���	�BI��^�P!����4�rG	|#F���2|p-�%��`�P�d�K��e����A`M����"z"�V�M�;����RQ���ϑ�7��Cr��c�#Č0�H5s��`�x��q��|ALjTc-dVj��Y\c�Vt���RR�e�å?��$-����bQf
s�)�|$��
Zg�q���N�g�lv�y?u�ɹ�����.`o*\�&���Pǃl��Y�ɛ���ʺ�����$�.d�[M`�Qd'�H��,mQev����&0����w����n�LhI�UT_U{R������5�b��"c itG&�`�k|��"q�eb�`@)
vF(T�)6�J�A������l�W�U��n ��C�Y �
���/;�*[�n-��a�@��w%X�li���G���~��XL�Ģ?��y�S���Vg2X��q0�Ɉ������GLV߶x��J����"빃��"�b0m���ii����d&����lh���m����E���>�t�Ͽ��Oa2͸D�^��d�#2d��.� N�\L���yxľ:��ŤJ��L�v� �YRӮ��Nd�M��(]Z��fa�!����^���)���Q���|���9�g{�\�W�.D]Ê�K��u<\�0}��	zVڞ®	��� �j��^�A8��n颤.����{���&�^?+� �`%A|<'�;rZO��C'(�A�VͲh
�E��F������~z(�B`�0M�<�O-1{b���?*�'Y��T~jNY��L	�I���|��e����z3���(�6#�&�0k�����aZ^����{Z�v�k%$�XV���i?[͛���?Lm'� H�!��M�i�+�Zq����C� �L�=kD$
N�VX�2؅��\6W+��c$H�e�3T9�8�,8?7	��3��m
�ɗjoH���^V��?4������#e��ſ]f��^�S��Li2�鼯xK�Y�-�Z��rA#d�̐qVܙ�Y�B���K>��чn*t��M�x�
��`k�u�Wj���Bk.����i�+�c.���6�]��n�7�N��.{����9�k/f�����Z+f��N���j�$�OÖ��)!N��m�
��֖�=�;�'J''E�D�q���Aty��Ϟ�5�{���� \Źw9�j�vՁ�`ϡ���8I�4�.�."gl/D�w��C ���4�l�-%?:�F��	;��f'�V6AU� �����B�wC�R����QOa���;�������q�P	_O��G*��\U���c��\�4G�x���fF�*�I!�REKe���2�d�>Zj^?2�u�gG�%uG5�u3�B�=F�K�Bz�Z?贈���j4�[{{��}J�jߥCȗn�8��z�zYC����!�Z�.��;-2�q�\��fi�Ӫ/�ZlEK3m�f�x�,�2 ޔB?��!��: G�2�\�����p���4Q���ѥ��-��=��G�0�;NGpt�-*B��\�9-�yKbaq�Dh��
��Y#Ss{�q&^3��� ��)��h����&s�g�I����dl�gn�ȇ��0V�N+X ?��2\7bK�lGS��(>����Q<�|!���\�@^XA�T��ꍢ��;x�3���2�蝋��IWG����&t&�~�`���5��"�xx��ڷ;�c��O>�#t��@u�4շs�� J�!��OIQE�闥q����^����>;?���a����.�L(�����^�S��\�g�6��Ώ��jE3� P� edL�y.E�',�&0�A��""l��d�LƿÏ��C�Ȭ�jKW����֗���f
���$�Z�,T.��J��;�����t-�A�R�kT#���o՟�j�7U�n��P�QՓ��ov=wk��;�u��cUG�m��}�X�,�+����@Ԗ���EUp����p�4t\dԓ��*:��"�(iد���
~&�8��h��A�����A��×c^zN
<}�f'�X�AUdM����ǉ�Չ�S����	*�}Yl�����-����c�*���!^�Y��O)�>k��.��7��@�+�W���r�[Z(y$ ���;X���y�X��#�C�K�#bQ��1�
6ݸ�; g�ۙ�֜p��.��Xf�E*	cvYIY	y�B�A�^�����S�g`[S�`�H�0%����I����S�sK�ZS_M*��*��oh��s���<�G��0\=�;i`��^H�[r/��7'S�t���X�} ���b~F;�e�j�e0����<R��6SS�(G�0@)IW���è%H��ۯ��h�E��',l��މ�em��hLC�� �%�k��SZ����"n���k�Dip#��,��������Θ�f<p>�#�l��;>�;��	�nfr��*F�UW�|�\���C�s�����c{�M���V� EK�� @� ���#��=9)6T3*B��ߔP*o��l�⪶h���q��- O�����A����*$&Քi�f� 7݈�Rj(��D��f��*�v��S�A�P�ۂR�F��-*AM!Un���v4s5�|�`��1[ǂ���'�a�S%���:�G\dB����!���u�2���� k�:%�4z"~���>��Tg�`��*moiIW����[FC���i@�\�N��a����*�[�?l��-f���L�o��K�v�bʆP��:�j�z� 1h	��`��]X�����B|�v�5!�K����
RWg+�<�1�ڃnѳ�~��c\�`��3�rG�	�#`kܪ~m��E����~��"��S�Z7pj�}ܤ�a�r������x[.�$|o��4-Lt��\�Y��1��]�BC���~֨���\�nkg#�w�r|�+�*ĺ�>鉼byL^��k�e�9a���N�z��dKdFޅ�-�O=��ӫ�»x�MO�1N�:�U2neڦ�je�u��{_��>�8����e�c�[%�s�J�rzli`�*^W��̳�
|ra��iˀ>�^5Cl
��C�X��c�pCf���=n�����C ��ި�lJ�[�alIXb!K@��
�&�+�T�L+�,Ѝ0� ���E7D�x��]�L���u�vZ�
�θ���Cď4��7�؋��Lkx���� �zu��%�rJDGs�2Y��J9'T w��v͊↱�I���#�~=�##<U���I��Zժ�;CFR5m�$�]�ӭǒ���<�� 9ؒ���b�~��R�O�+9���v)�wR��Ge�������$�
x+2&�"�ө���F(3\;6-���:8�N:��c(T�2�����4pU5>������i��INq���ޓ��D\�0 �̥Z�B�<�zxQ�q��+ʓ4qV03�	�)3�2�C��j���Dרo�ƿ_�0,���ȺX�[7OQz��A=G��Lg/����3�] *�5&V,��\��)�qL���X]���8�ҹ�hK�'B{*!�U��%wiI�!�2��I�ׂl}��u/����wN���YW�N!��3*�#��)�H(�[v,�e���OnW��# ��4�w�H��Z�F���X����Q pD�G�_QD'r](8HTIbz;;��I1c�7�ٜC?��&��~!*�t��N�|+�5ѓ��2:Lu��<2Cq#z�e�]�\�Y���:"�ԡ�-R�#ܿ*���wS1�7��O� �j�Q��d��s�m�']MC�E���'�I<���]���\���-��^�I��S"F�s֩bS��p�c���R����
�D�����K�PF��F���IE8f�Yc+���W�:{4���d��4�Y�b�?�~�$�u��y/6�4�RF1�����ߢZ�����v�#��D�[|զ���)��L#�~d��~��S0�/^��j��.�s�+ܞ)��Z� i�a�"��S�vl�� ��96�C������q	����Dv]f�����ӂ�:ǄIw��-Јݏ}��IpԿ�x��i�b�o���v�vG��8l����}1v#헃�6���|�+��	�+��&�D�{!AY�T� +�js���x��F��^{ٍ�p[�WTǍOK}2�,K�I��(�O�>D��B ��>q詘DO�1�޸�
2���ď��f������D��b�<ik��f: �Z_��*P�l,z��Q���c ��ؒL0�r��.�U#��8�沐Z#
�%��!��j�+�d�&��r�|XE��?��$�&��Ӿ��R9� ��\���ӿI����~X3g;�|jJX`�$�}�C�(*�(��KnC$�C:&�c=1���~͓qa���TUb[�a�I������	K��+�\��(!���z?����ʹ1�������s�>�	�l�ËM��6v��8|�L�)z��b�Y�� ��J���Ik�u�!%����C�Pq����V�L�
�f��ǧ�A(�r�ܢ��B�P�|��%lZU����q.�[���f;��g�ن��(>Jɒ��O~���՜��2	�������{m��+�ܜ��i��ID����&�B_�$�e��?[�e����ԍ���C�3OGf�KN2�/`�"4+T�;��Д�_ �3J���ҭΰ���y�yǻ{b�����5~.#��xJ#���@mg}?=���n
��h�Uh��t��!]������52�5F���tN�K��+��'��Gq���S͘�؛Z�^�^ǁ��#��n��4����x�/k��d���~����ł�L��
�� 8��5�w��% IsXƚ2�2�@4I5�θ�s���������.���%쑑�v��%�%1��r�dy
֕7!4ǜ���DN6��}���?[���3LU��z��<�>P�
_D�#�������'(eW�O�虊.#}	��V�;%q�EmM���.�v��y��DA��:l_p@O��ǲт��.j�G9��xN��|�>o@�Aoz�>��=*Z��Cnj��e�Dw��#��\ǘ��t�|:�L/%�F����������38d�����k4ǲ�(C[?ܰ��:jё/I���PE�6�k��{�*qUP��X4�r�w	p�� ��K>��-�)����N�n�Q<�������q�ђ)�s���DqU֖�b
�Z�S06Ă>ʺ�r�}'nl8_��Y��@>�a\�� ����{��0i����{$����m\��jt���̓�^�|ո�w�&{5J.�-�*DP���C`�cők��W���k�ֳS�R~?p�9I�w$��h�3_͒��
A؁�|.�*�>8'������bZ���$Wƍ|��͸S�����D��xo1B<=\�*�Cv�v7�r���X೷}���Yq�e.5��h�7����R�Ў���P���,9���I��,�i� �����lGY�?tD�(�M�O�(�s�/SMP:Xbu��+Yz��_��W��}�0 r9�7��1���-_5���J\�3i1�9�d�L��
3P:�t��E���3���a-|�|��Z�� �����<@Cϴ⡁F�p��{�G^��R�rz���	/�֑�*�mjAfQHVZ�&�K^B�%7�w(�.�5��X	�=�i��p﹦��f���ǈM��_I��ųC�����,��EhN�lÁ�Y�,w����R� z­�$�k�l�.aXZ
TCJo�{f����-���b�6����9VYz�G�r~�ZxW����y_���gOd��2.��esDЋ9��%e�oxK(A��?�mm���b�����TDϭ�z��t�(������Ŕ��z����\1�w�`Ѡ��l[�í�nɾ���H�t��A��X�S�3��׏�꿅/UՓ�S�������f1�=�C����V�$��{n�Al��a����Դ,�K�d����ff��Zmbb�}��u�R�4j�Q�_:mʁ�Otw��/}�]>����p�"a��5e@��j6�K�Gb��N�h���Sx�-�x�t�i�z���?�IzI�p
xq�-{c{�Ǫ�]����2����K��_�~�~��U��-��gU��\
mn�B�ob�Z�T�ً�����a�v=a����ͯgc:3�`�؂cp�U�i�TGF�����d�tx�����-R�
^.g��CQ(����'[��xrx�
���'"1
�t����f�J�{?_��78a�*&�����b4��D�E%|1����c={�2\�����7�sf7�W&{��3"`Grb[�,�X��$�}�����wC	��{�A�z��������L�iBondڢ�(�l<:�Xm�O �@Xr��@�>X����r�
���",�X�/�qRC���Y���1��T	�M�"�b{�n`=�v�Z�>��eXwa	��u���2h���E��.+�ÐE�{[�|��xM,�^�(P�)� &��K	��L\���b!K��B��O�rZJ�F�m�ڮ�J��� �B=����_����i ��Cz�E"h���q�Wy����;�ݠ�\#��	�W�rp	4L�?��p�t`�iP�u�ݎ�}��D���t��a�!�?�{�Q�rǏ<���t��}�G��8�yJ��#�{|��_��{k
<TC,(���Tj��~��e�1M�:;�5i}�O�HFH"?~)��J��ء���Aʻ�����K<����9i
�φ��u������2�� ZD�9�5n���BƆ���oϑ���8 !�"��A��J�QWkܟ����k�&t�$����B�-&���9��k�x/��4�� �����s�Ԃl��>3�[�:!]���TT�;���2E�)r&�H;<B7_=�&����K�����f%c1d������h�Su��Ӻi`y���P��g��4��dV2ז-�c���|�3B5�W�gO4�%E�e�Sb��X��9�ޘ�'�9;�[�+nq�e����Ր(c��z]W��vR'P����� �ֿ�t�N0�����t�A��Ie�[D�4�9��Uw�5��"6e��9����^�o��0|˜�RoV������S��e��-G��rQ���x�%s굯���֖��&�T�ɴB�.�5��Bf׀)"dVF�{��i9�Wt;��*�a˵�"��&bW�m��u�C�O��@M�s�
���d���;R�ޕ,�����#�ɣNW��[H���l�)�MWM�~WHI4�E_��1��\�;'�p��{ִ��H��M�T�p>Ӧ*���p��i��uDB]}��Gm�X�e�f���P'�~5@�c�hn׼��>?kf��,�I��1�'��3�U�|���}�K�`���1n�-�v�м�b��~�����I۞�V�~!�ܒJ=��/�V�(�A��h�����I�C� ��� W�j�{�qz����;OO&�|�x�Y�:�Dty��[դ��ޘ�&)xNEk~�a�ѩl��BRg�;<��H*ʸ�C\��DR*݁�WN&� �\��=������a����?H&�I���էޞ����~����{k�c�����Y|�yv#���G�nWD��R���U�A��M��0�CK 4˗�?5�W��B���DJ�c�,�h�=��j
��/fL��x�EŊ��o/ Ա*ι7��u���i�>Z�\Th\�_OJ�$��qm �#S���?��X����ǲ��sM��9��:�G!�y�Y�6�)#	ԧ�G��~(�h�ܪ�IE0���݄�Ὦ˷:�8�U���u��ys��#O���Y��ʟ/���զ%P�Aq�2s/�d#L�����,��������V�'�Z���ޞ�*��}N �Wߟ&j-è՜�Q)�;�ҡ9�7z��3%�X���lYHF��&e�ݧ^un������Ә��o�(�V��G8�/��e>d\�X����P�О�� ��v�����4�z���r�q�̡��Vk�;�v"�rc<�P��?�nC�L5��mh'��,�%� Ѧf9�F\g�kV���P������1��O�=+����HW��"'��`U��YS�jo��n�
g�&����W!�+/5;�%�c��s�$�V��cO�@/%��ؐm�8oB6R���NX���~�SV|�GmȀ@$�[up�Tz������2IV�N�٩�Ԭ�=w�*��g�E�AP�&�����0���v�#�kY� v̒���ɻ�"�9]�82I�V�J`'��ָ����0dG �����g�P�}���`��]i����˲!��3�[KhbQq���]%s2W	`)���{���r�y��fk�$R�?sc�^~ vVS���Й9�}�=����4�AoFh�礳��y���T3�!��D`��b$7C*ώ�X��2������#�+��EW����o��֋!�_Db��I�G��\���H}���!)���G�A�;*�� x�Xp�2��n�y���>����8ز� �^���I���K,v����`8��C��a�ᾴ��R|��V�1��X5f|�L�v(l��dMA%�W��ky�[��h �pO�{�,��a��j��_��і�6�=�u�W�)I�Z/<jb�f�4�n�:C,��*�c�����狮�-WB�ʜ��&m���L�yJ |�F�A��!��|u_\T�A��[���9Ii���uG1<uk�����ΝS�;��v
��cS	���� �;��E{�-�,���/+�Y!|��b��V0�4I�	�t,�*���s ���[�|�N���v�4/a՘	�=8���/���8��8k"e��A{�U�/x6�C�L��=4HP��h��S��)�J@i��x��k�y�@{@�=vLU�D��=�{�TX?K� �����v:���"ιeX�U�ӊ��̑FW~:��V��U$J�����w4`1�G�x&�o;���'i17�e�>i���ҟY��g�Pmb�:���n>�zi�^�2"�&��p�`N�$g�~����(���\ݩ�p����+%Iw�K��� crWys�h����X�|J����t�z�~qk�B��p �R�ch�qb�^l:�i���z�x_3�[e��6O���N���Ϙj��XTP���|���О�^���T��wR�=3���Ű�F/?t��`��>�͂"8M�k�&����4��O�_~�����dY
�b`��d�ZZb-�ݾ�'��s�n1�����C�IUoĿ��rn�W�qZK�R�ݣC���(��]H"�^�Hb�U�Y)O�T�ё�s���ۼ�6��M/�﨑����ߠ��'y��mG_E��Iݗ�/:ani��c[�N�\O�ޔY���5��ރ�b��a��S�;��I"������A�"@%��i��=A\���wa�(���gc,F��w���D��O�-(�=1w���,C�-����u�Ag'�k"������CE*��+�#��w�$A���v��R޺�i�t]P�o��O����1������D�Q�'��k�!�q�Y���׻ӑ$��AY#�"����A`+zi\����v� ���kV,�GC����[�$%�m^�8?}���b��!#��d#B�o��-�L�����% �y[H�Z[4��V�E�?�z�/���80���\�Қ�=� �6���0���>p�u�d'������l��H��)�M���C���$�8IW�U�6ݘ��J�nU����?�G�w��6Q�?#���6���&G���$u�P��Uu�켊L�,8�cq��������W2��AF� �x���˝�|i�	1Ɉ�0�֕����: �]�S����I䜩ú��x�FV��3�����
��+����c�|T�J�<��뜤�B�ٖ���e�j
whb�`�~��6�Ml.�O]����DDU���p�&�.��G�O=������4�cR��ܬ�����dY�ܚ��JS2Eu;�+	2΍��4�A/���G��k���`��[o��L(��⓷ ��j����cpb�i2KO77s�����y�D�'�"�������4�r���|�R(��a%I�ˉ(�6V������ �/W.�r�!DõZ2c˺�mA�*
����_�sN.Λ笃ХɉB�ŔnAU�"��[g�<I����O�k����gכ����[>E������
<u�[�����z�Ԯ�[1ӓ�}�ǂ��gA��RG��J�ᚓ�j�M}Ӓ0nJ��ޝ}��h�Ș��Ȏ����� ���ڀ̒.�)�YN�p<y:��M��!h�5�g�7M�E�6�ޙ<G�,��L�җ��#����:�]��Ë'	�&g�)��A���Sĵ ��T� ��d,�Ф�[tFfm�A�B�x)�������J����lq֛�G������E:X�[>�`��i9�@eХ\�{LQ(<�IFOz���sD)�[z5�^�2�!+ş���u%.eR���ܤ�?Hc;\`����?�i���bP��U�ps.�6X�� ��}g�F��V1]k��TpiXA,^�M��"X8���`��ڳ��B�_�<t�&��P�u���t[��E�{��q)}�����7e3��^@��Թ���e>�Ni��-��$N&�G�K�^��=���~{˩8;�Ӳ���\9���l��w	DM�{dwqEI���j3��ߨ��'������N�S�4)���������j��p�TN4�5 M�x��ODw�Q���Y$|S3t�S�?�Y|�;���ۮk�3 �}�2z�q[��[BS��9�����f�2��i�d��m��"��'�.�L��Ѣ���HC2�2"9�`fE���ùV#4߱��f\� vG�=����p�A���0��oۼ�V &����d���������p{�oն���i��y�	H �% ~*��%*�(b/&�Y��NQI�i&�����I9Ϩs�% ÿh�^a\�a���0����~v�K��Ȍb�1�g�i��چ̴�5l�GS똯o���ӧ���L�$�Q�������)�n�R&���s�V<����^���[�l6\���[�0��e7	��Z�3JD8��'pܚ|�PkT���JsF�t��⬭��e�&�s!D`|
�	���D�_��A9L��A�¶<�@�Ix�mO���Ĝx�<t�����/�Rc�,�S�7j!�v$�L�r$&�7��؋Q�w"C^/#<,�A�J�w�6D�I�h��a���!��q`~"Q�Gp��R�\�v�އ]����DCd�������nUj�^��:8^��;*JjT�5��En���>���^_(��R�Jm�����hge�g@6��q���%�V��e��N�������+jѿCc��3��U/&e��P���G	��8�Ik���V������WT�Y5`\����w&��I����o�	0�/z��bJ�eA��tP�����!�=�����y!P@��px�QHU�����r!N�NzY$�ek!1n�O�^�n/eÂ�b�)\�� ����_�Qv�;UB�5%my=UШ1f3��/���=^��L�B�#B7���$�� R<���!B[7�"�ϙ��"��4��.j�[���D�|��p����OK�pĜ-j���cs*ֳ�>�@&��ix�4*�Q�P��n^�4n��X~ъػ@hJOÁi�'��'�K�m�ES�⨨��k��K9�DXE+����nA��&<���0�
3v�:O�p+�#</X�������s���|�����zs\�D]���a�Ci�tS1��z�P/�v�����D^� >�%*PS��qx.^�,��:q�&a�
*^C�t�a �Zb@ڊ%�qVR%ܘ��1�$����k���7�R�P���)�?�� 6�G֝�;�=�f��h��n�J���`�|
u�ʔ�>��rA����B�S�~��]ι�y�F���c�u��g�WU����$�4 1�h�?Ǩ�z6���a��ߊةq�r����sXqg7c�V+�Y	�#L�&ę�@�	9Ga};�2B���x����$���`�}��W�KQ�uK��.\;���Vk�E�эwc����_] ��yv#��$�Rj�BV4���C�Y:b^Ւ�6ω:�i�߁������8�ӣs��I
&>�k���CO���������u5�z�(���?'����JX!D��c�}��u�%,�T����z2�0�cw�'���`I&���q'�D����d���].k�[�$a�:��d��[j3��(h]Q���:���kȒ�:#���ހ�g����
?(��?)6�uF+�r4-4�S���,�S�ǘ��˚����˙�?�BT�~}���4�K��1�t���3f���js�Qu_S�#���U+�d�DXt���dD�����&��A}�N�)y.unU�N�	����nğ�Z\��ߠ3���&��:�?z	�պ~�[m��u�N+.���Q��`�2!�z��菜�Q�q��,��0T���9�p�/V�c�=f����*[	ES���^Œ��a����(����T��NJ�XD{�Ƣ�4��s� w��~Um�Y�V�.fV��%�mA�g�.��ƴ��nχD_�u,���*�GK���1ˁS�
�^x|�iD=�:J����*�u�K��/`ُM;�29W�ж�i������<�ae���=��'��Kq,��ˁGx�O�2��z��w����.��9�����a�	�Ӎ��m�"H|��kN����FW� �ī��ͱ~����|��N�Э.����v�׷��ڐ{Ҥ�1��U������ǜx^�1_�B,���֣{_�Yݛ��ˋ�B�6I�N%s�t-����0��S6�	���S�S
~Z������rR�7�B�a�!5>��XQh4�wk��U�KŨ�VT�	I���'���o�5��A����kq�B���^�������rNQn�vǲ�}� �=&V�8��e!�q)j|����qK�j��I�"y��H'�
C4��Y-����)�c�l>z���6Y�}��k�R�}�A�WL�_�,���H��f��qC�{�QR�b�]�]G�������1�L�B�'=�P]�Y*�oof2-J��>׃';�A����TNr��v��P�'��1����z�� �!v>�0��SH��J�=�8Q&�>B�D��>��Kv?[8�F]
�V4Z��=M�zS�	a�~�r(~�o�l���W����dR�te8�^q���3�������ڙQ-3����Fe��_Ķ&�e����['�G�+d�c��}�?�)%psN 0s������]N6��&Zí���{�Yꧏ�E�L�_�s��y�(���6S9��)~xz`���(+]�!~�9Z�[L�g�ǎ]y��✼�����b
�f�x}U蔔CL��*Nj��{�d��h	���ޥ�Ƅ�h�C��+D����/�C%���w�K���z����_E�<��!�R+�M\����A5R�b3�5Il�y~.2�h����,�޿��ե�8~�e�jȕ��ȃyyR��.�`�N�Y�a���#r��rI4��D⵳8ޙ1�8��!�1~��s�QN��7Ě�<�S�bĴsqC��N���΢?c�sWǿ�:U߉�M(�mөכ�1p��R����O��e�j�n�]�^>�֕��^u�a��*�+eY��sn�Y��gh�	�X !P-'���)�N"`�K�D�*�v��
��kb 2G5m|㼔h!޳��k�3b����(�K?	[��AĹE�Ҧsu(�M�n�9�{�L1mf�(��{P�Q��Q1��%�c���WTq�T4Ǹ<Ze9�o�"D�T����lEF"����(E~p.US:}�S�� Q�[D��uΧ��X'U��ɽfc��t����̱oȾ[1��O�l/UDN�/�����y���f	8
S����?C}F`�?��U�'�Ǡ���L����a:����J;y�P�9�$w��.��!�+�l�V��mE�E�ܑ��YJ��+�<����p-U�i���:�̶D���Ŧ}�)�Bs� ����֬J@~����|�{3n�(F��'��cq��G{M5?}�jF'tͲ�x���+[�)ȐG�W����|mn@9�,���V��C�E�M�����H�,�XPj��j\���}B��}$���bDh���#�)�n6AS��1猙�3��X�=筈f%+3u}����uf���Wa��+��)ۛ)�%�8R&�_qt��v�l����~pdD��t�[������%�k8�l��07�Q�ް����\]��⤐W#S4�t�du7�^�%��ڡ�y�O0�Kr\1Y��*3v��l��5�G$����Ųإ��}����-R"�9��rq��e�F3)F�^׵���e���?z�Np<�.j�U3�؝�v)o��" �/R��&�[��*�3�:��W�-��M��9���9¢ё�N`��-Q��tgX���3����M��6֩�sk�8*U��4�b�M�i�u��JW�% K����V©(ԓ�?Ăܱ�AUO�$�ס�X(J*�X���zm��YRk\�p �qp� �a������;"~ś��=JEY?�8
��v�ӈ�P8R�K���Ӧ6�u������`RQgyVV]v���?��:���@���1�� 1:'�nٲН;/)��W�%�m��⯢g/2D1���'
4�>�}��f���|ܥn�ҕ�cg����?H�U� %��@ڹe[�<T���@xL�:��=pl�^ʏ& �.*\��πy�#\Á�EM����.��}�@*1�X�z]b������਽����� ŃY�C�fb���,4i�������������`�cM/��8�9eCQɘ����9����'�\�� �R���)�|ͽݸ�cb=U�6�M��<N�{,'(�+\�ݟ���ѩnH�F�Pw�}N�v�S�{���z�4�uC8�y�G����܊��"N�3�v�O�'YHj?�΀�`��MB�j���
��O�PzKt, ۙm_;�y!�pR�)<�j�5����	����#F"E����(D|R:�����7QsQ.�h�o�En4�	�l)���ŜV��<��u¶�wI|w�N[�a<������U�f'�-�Rg�5�ʃQ��C9�C̈^�]�h7��=A�6�;P�B�չ=@uWO2���L���U����VA�5�a�R�(]]�? �Є���u��o�6?Z��N���{�2�}�Wdo�L.m�^���=����z�ݾl|���}(e�~0:pW
(��B�3f�V'&�ޥ灙��0�ܒ����?���\NZ7y��S�GM5��ل���uj��z��n/�񵅪
!*b|Fb!_=g<Eoo`��hZr]��t�Ab� "*�Ey� �䒿w�[Y�ԣs��5T�S	Ŗ�3�{��`V6�����' nr]j�p�o)��|��C� ӲT���%F����c-�L8R�a���)P�(�7HeV^D�J�O	O�<	*���/"<�9����m�J��:�w��9�Y24=jmXBY�UB�_�0Zf_D;vt��P�� #Xu�\aDz}8ީF�H��z���͏߀@�7x���
�ۈ��Ň��/��fic��o�ӥr�n���%������8�V��!A��=���NB�8�WTD�����C@�K���ý�����(MZrf�}�
#TC��-�
س]���=4>KH���Ն� _ɨ����pZ��Wh��2F�x
e��y�N��e���z�o9�I��O?dOkA��-BbQF%�4��տƽs�gF`nhq��L�׻������3�6� %3䖶��E���/V��6
���)����-	���ǯB�0���%m�#�x�O��!?w;���(KQ��W��#vf�#��ZTI�����4�7���է$`ֈp� �&����Ke?n�n,����(�� ���Y���Ae����V�e��fD�=Y��y�ǅ�=ܦ���j����N�P:�ߎ�u#�L?Õ1M�K+z�۽O	B;��cZ]D�"ZQHc	z�Ӓ}DO�js:t���~dD8�!�|QSB�����T*{YMwq�z�ڶD�N�h�/jl�(�'�H���>'�;k�J����_��Gj=3�4�1�*X(.���N�r{ޅ��C")T���|H�m�EE�Xƒ����*
�,�
,XU!6�/+�^4�h�R�-�D���B��q*L-p���>�4���R�Ժ��N����z�� m�b���4wa��а�#��U�4o���
�H�H�=����f�6��^ǖ�D�!�{m��U�j�D����t�C��M��*�g熄�%,��8��H���}�ę�>a�
X��)_Il���H���� �K&�<Zi+3�7�'?��m��h
��40Q�&�z����X��(Eaz�3W���P�����T "ߍ��p��Y���L'��6�&��d��;��R�Ȥ#ȱԪi
5�S$T��t��|�<��PR� Ae��cŕ�n�!���zԭП�h6y_\
�W�mUqz�k9<�3y���1g��f_����6� �]#�2N�O�z$ֹ�grmm�O;�H��	%9I������r�sƒ�0�E�]m�l�bQ
�����q��q,v.��cL���G�ub/��:�(1iH��!`u�$��������#��I�K
�cimBc��c�}0��-P�qg,���%To�0��d��r���'�S@*�CI%2m��K�b��_�/���]I��D�q|\��%j�MLYFbXmp�e�2KH��S�����u	N�3�0ڄKe���#&���<�_�=�cT��G�i
ߧJ�G����]o+?ݽ9%���]ɸ��� *� Ǣ(���˶]ZC�iӀ1h���|Y��0�ƥ�7{����2�����, 5�d����~͘"�T�&\�ݠ�ז_{s�g��&]J���*�{�<����{ܰ!�@��XJ