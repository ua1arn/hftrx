��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY���Q��3���Ss��t3�ɫ��zzm-!��#^�g{����Q�LC�k#��q����
w�i���]�k����X��Q#���U�[��åV�C�E[̘�� 
ݼ���T�.1Ҩ;�]��`�Y
��B�b���UhZ
bRH�1:�V�%
���Z�h^�}��۬���fG���0�B�a��F��fA&�m������è[�Y��g��2z���p�)ȥ���F��"M�x���M�}�j���R,�j&��V���� ��)���z�;�d���T�}���}{p�x��+ۈnq +�d��?~��@���I��g�����e����r� Ն��K5e�L@�(E!^4 z�n�Нx5��Tnu��EdW|��*}�w�S+ע��u(�F�61����I"B�g��cW��I|��ـÖS�v+�� `r0:x#�81[�T�Ρ�a��iX����jk�{��l"�xGp�A�)�7�c���J|�a꿮E�
�mJ�]�L�i3�Ӱ{��Ǿ�a�)� αKHh�. w�7���R54�;��A�ؠ�,�bT����9�L����0Q�*�B�P{e=B�A��G���w�]]�s]�d��_�H�+Ͱ��ݘ�c��,(D���t�A^RhG�Wz����u��5��P�m�����y,��$ϟ�އT�W;l�2 �;����!K.�Z�Q>%÷Ǭ�u�Hӈ(eEɮvq�ZN�Xg��C6�z�!{�C��U���J��V��S�ሁ娉Q,&U�%�_�<���J�ȇu�Dl�%��u01-9���g_T���%Mq=7�wD�3���&���A�=������]��DSU�a�T�@�%3�ռ]r�4gB� %�n��WI֒ႋ�N��6�r�5�;�Q߰�T�߀�Aׯ��,V/�I�A\))� w1|�iHv��Wq`k���/֨�f�J��uW]���PS^?6��jh)�6���^���9%�S��(1�Z�k-���.�Z��S�2�uF5o<C_��*쏔Jm�N��\p"<}caQ��]�$ڦ!�|=����jE�Q�8�S�Cm�~�Z��X��i:-�/`YX0o���p��?��-�$��_G"�ϴ�sC}���	���j���	B��%V�#u�?"��_ne��)>�ܓ�k�������Y����#�ctq&N83�ϴ|l�w�=���&�50Fܘ֣��~<�g���i��e���ͅ&�f�ic��F#�ר�ʤ�厴��u{��{�=�|�n�����iW)�/Eҿ�t��C�3����a���L�����;ה��U�{�{B�|ejr�8hB}c?���M���=S�<SH�L�%rc@�)𻀳��V
?����bZ����=H�	�t��}�]�x.�ɵz��:��.F�Vd��j#,c�u�;�Y����|��&�0������0ԏuwP�0s}P����/m�bұA?_R��{��C���7n�҅S��x��Ap�Y�(l��c���#Gv��ް͎n�g)$��EZ���YF�c����Q� �����|�M�J�5�T��3���Xg�Ūc�C�_�3�E�����^�@֍�Vޞ��>#���+�O7��5#�<�vr�G>\�]���F˶���-�.	1�ܝWq[��g0}��ٰ�r�;7Y������t�aX8��FX<%z��12:k���IC�0�98+���q����S5y�1�Y�d���S*jUz�zK6(_D�&)����Y�X����s��o�s]��hyY	}?d��[z�V*��}�^�0����Mf����V�A�z>B)\��|�XKR6եs�uD�.5/�0��s����c���1��ʽ����H�
�we��	��5x&� �s�R2Ӵ�3�QT� :�,3��I�<��'�b����1P���I����H��powf�� ��3��wC�`�V��F�9��*�j�|)�0Y|�w�%zcK;�E���Q�ci�+J�o?�������+����Ǿ���xt��WJ�nN�y
��=�>�6�:)qh�ys�G}�_%�}�6�kZ�h��Q�$�ՠ�͞+�R��8kK�����5Q���<~^H=*iH�Q�X�r�o����� #y�9|�)k����˩y��4'��$Y��f0H���BN���P���Di�D�B\���z��.�� ��Ֆy
n��	V�mqv�Tv�-M]1u,�*H<��f�dJN$��ж��E�0����}�m�߮LW��q"G�`v [�bFu�D=�S��&JF.ە���t?�����M��������,&Q�:�:��f)N	��BH�z �6������LS��l�e���R#9��hr7�j��Y
A֌R�&���B��*���~�[��6��
��k�C�T>X�a-9�r�qKYs�i=���^�8�mx��T.���?��2�QC��ba/��z�������kp����`[C�*?U���䳃��A'#1��J�u��h�>��d5rM�;�s r���b�OY ��tָhL�_��xd��}�S�E��rva�aS���V��9j �D?�ԥ
����]�e{���$g�k0�e��6z�689֮q���E]��=ظ��v����%!N������s�
�=:&8{*�����=D�=K�iUu���ۊ�Jʹ�p����͗�!�D��׹�fv��J�BR�D��u���0�d�9wd�s�YO��br��?���|R�:�W�Iۤ�$G{>�vH���)͑�as�"s�u�M�O��/�C,S�1����c�|��Z�b_�z�Y�y�i��-�31]�l��NM����h4�����˓e8�D5LI6�x����