��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`|w�1�����%���C+.:t��v~0�dtH����Uz������K4�w��&��'o1~)���6D<�RbvZ�r%����y�E�i!~����<=�ә�ⱟ���1(C_D�-e�r�����&u�&�L���;�4�.��Y��70N*,�a��Bx[�G{���4�]m*ɻ;Ȫ�
Q������ӷ�Jp�)���1!��py+������������Z���Z�ڰ���/��� �I�݋�B��j�ZP_Md#W`⋙x}8fBg���l�:�P����IT�L�r߫�u���wv^���Ir̩H;��[��R��5����M[y^A�$��nݾ&=��g��� 5"��^s�1�v[�Ũ��#Vr��S?�6�4Q�\��D�n�����Q��,���C<���Oƿ�&uk
��X���K��$�W1��|*S��,��`��<�tKh�������KԤU�N:_���^�~�!O�4"<�6�R��:�_وj�S���s�?��d�'�vT2�ŀ0x4��'�p(�+����f�E)Si:�e����X�I`�+�p�x8�AS��|u8���&�v��+� sQx0��"[�UϨ`�j}ٔ/?�&�&���YzI��M��Ӝ��6)�L�
a�q=*�5��4�%�5	�gC+�mb[�]�������ʉ��&������C#2�G���{�
�tn̄^���Kh��q�[�3�=U��;�g����rՐ��/�u
�$IY��ݰ�d�n�tOTYZ��R�����G�.?�;��sS�Iꫵľ �g��l�O�����qT���W�3�?T�>��ؘc��;@ `�k�	'a�]�ɱ���.{�!��vO�v,8FP;�<�ϩ�_��Z���<�@����:Κ����t �oK�c*������s����T�˯tŻqu�I�QoK��ь���X4c���ÒZ9j���-`�F����}\9P({P�2�6f���H��^Ga�>Aq]Иt��u��.)J+f��on�~@�/T@2t�M@�ڹ� R�ől���ܬ�r�d��w�܉�	|uXaU������嬯l�H]$��0,��=\Iŷ'@գy2 v�.���=�A�:,�# /�pO4�{O��� �Q������	�?=Q�%� E�B��pɗ�(���a�5��`���M�+ g#lh��G��]�R
��룑�m$�5�}�cd�Y��J�	�>�sk1i-�G�I�D�e⨐����Y.�+�ě$:�cc��#6n��$6��e&�
�t���n�n��|�g��f�W��)�$����x�6�0�$�m���9n#?�!bmy�VEf�c)9�o	�� s�e��g��� ��H^H��6ĥ�A.3�^�:D|[F���D�� $���'o�S���'�`�}�«�1C71w���`Rk^e�͸���]~E�/,��������F4��M<�R�g�%^�a�}�zy?��z��-|�4�m���h$|^��槇�d��	 �J���� �y���` T*J&�z�ތGF�%=�p�r���#^<}4l|���nQ"�	C���n��fρYbBN�!F򻵙���ŏ]U�͢b�	շ=�&Q�m	��w!�����5�.�F�o���枍ft�C�ߜ��oY�ʈ��b6���:I�k)����8,N�{� 4�rx+�9���NiԳ��"��?4��|��<W�6�[�
��n��pR��\.V�4R+F5��b�㗔vu/m����Glp�؄�U�c&ޜ�3eC�T�;D��p�1hm��#t����o&�����ڽ�v/�o���/�H����S�B����a��^�ҭ�6+ ��q��k����UH�"�qV�w+3��_7|�z�.���1V&(vj_�G}��o��۰��|�[�9��}q�C����V曧����g��>,��+���h��{��iۆ�����qJT�)�*}�5U�R���B��lx<HV�SNP�ə Ύ�������ﲽ~�qB��5�Dw[�F�?7S4��~� ?6��T�E��&G��L�CS�`Fͱ#�ɸaw4�Ϣ�����?�˃`�(q����Es 8ac�q�Lnܔ��ɍ�v��m;�+�Y��5�MM0�(tK��3+1}��\�o���y�Gc����?Hk��j�����������9j��x����mV�#�]7��`��|�ꙋmMW4F�HtM�+ <���e9���vk��M��_V��F����-������i�*�^�|o����˶TLtp0�� s��j���{�h~i�7[q���M�����[��T0Uv�;�P�N�xIY���rh�h{�e�O�5Ǔ|� Μ�d4;忼�j�D��1a'�#nR��m�����ȋ�:�Y��(켓Hӛ�~���TAU;�T���p%��J@`;�I�<����W�����t;�c�������/�Xb�\�E������Ha��QE덢�A���%-
1����s�"��o�>^��A�_�R:.��ސ>��n4L��XE5��5�����;�JU/ֻ�	�K
�������xl���%Wժ̩ߡ�	�8]J/A����v���,��W���lS��3���s];�U�X!�̑	 �^��me|�ġXH1uf�G�z"��:t�L!�Q
R���_>����.�}�,��e>����"@�[S�Wq��lr�~��D3����̍	�@��թ�����o@Y�=z^gKh�䬑��bs�8�l�T~#K,���?�R�X��D]1�MQ+��+��zI����Z��o�W��< �|N���S����AH���i!�:�`����t_E�HJ��?WĨѰh��RiO����&}�*���B�l��o$�UD����Jm�QB�-����W�I���F�×}S�����#oF6~?O�~��~���0���t��>�[��a,�Y&�=TCK�ĊJ���X��.Ýx��=x��<إ�O$[ޜ(s�輕!+4���|��`�9��XmE#�C��r	����Z)� u��BT
��и�`��Ǆ��Ғ��VV5���A�!�5��P����sJ��vPb�f-���SVniGmE�⨎�����ׅPm��L���<;ҿ��(02HC_>�X�ʵr�ݨ&a���S�.O�e�g�B���M�Ȋ���n�^=�Q)�v7�MR#�˛��`ƽY�sL3���PZ� }|$G��n&yԡ����O����ܚH��^m�[�pQ����6�
v��E��Z{e��[�9e����t�����v��mj��ȿC�)��伏z��Z؇^��������Aslr�����X���i��_��'�x�a>�D]�ϘӢ0��$)z�� �5B����n3�o{ޑ��� ����V�A��i�/WY����h����C�X	�#����+�/m��C+8L��pg1��RQ�!���)�nϫ�r�&R���RK&�y�SKt�T��7�s�u��o��d�G�>Q)��Y�X7�Z�� ŕ��5����A՞����Jo�B�;f���u�����c�!�p�e�+9�#� _�9;�1C�� ���j��4�2��D/�׬6���˙$�[��g���Hn��J�[7�sքyg��?�cB'��Liae쯆U_��GRdH}z����1(aoY��O h�����	�'��V�xt}������ԡAR��Jbi�=|m|ϔ���$!!ãi��!O�ߘ��A�`�l)��!�����P���9�.�K@ǃ���#Y�_&��2pEY��l��/"j�dr���9��ʑ�i9<{-���*���K��0�џ�}��D��~ɩN����C*o�D�m�-���g^=���"���0��ͦ��2�Z<�:�
�[jQ=�����1T�=�H�ⓦ�h�(/��K]0�b,�<P����Z���F]��ewؙ�4�h/-I�ю���V$ݲ_U�:��P�O�z��W1�8�%	�i*�W6��X.�E����Y��� �����?a���� ��^���OS/�J�~7=�u���jF��
Kx��4����oNm�@IV&Fg��{ޣ�~��	U����ŘMg���*�g��Xʦ6p��{E,PK}�C.��7���g������cm.%p����e趴��Ŗ��N/�+l�-�����i��d������WF;��m&4������<�Y^��|�U�4Y=�ެ�x%�8]J�o^�c�ȝ�n�^ ����g�1.,���)��T� �͉x�|�x�>̊���sq�"���[1�a��RVލ��<��G�?J��1�G��LX��3^9E�~�Ζ�����|�Q��L�Mل�Ҷ�#�FJ	#�|�s�M�#dKfh�/U&��=}yUz���i4єU'�)�SVŴ��S�H�����x�"��������`���џ����S�T���h��x����
J-��l�杜 3�H�qe����_{k��n��'����k֮���"û��"Azn���]U?���NV}�.���2��#^ z�/�pu!���Plw�&^�&ư�@2c{��7N+��;��FW�.��2����֗�y�^�����#�v�Ae���-$�8�ﺞp��)�M
��Xσ.��Q���N��&�������/��$�}wT�p�vf��l��\�:�l����P�P$��k�iB��Ti���W-=@�y�4>��	L �#y�]�+�9w��O�6h�3��ki�7���l���ւϦ���\`Ԝͤ��"�� �t�$o;������!�)��/H�l���ǀțI�8Υ��17��j�/|�D	.$ߍh�I �((��١PN��	_�дO2�m�����I.e�
��7�i�;���l�����f&(����ǖ����<�L=�^Ȥ"������39���PT��������H�Vk9k��;�$q�WD���,�Tr�<�*k��w��z0�|=ìMA����#V	��m��� �66�P�sٺ��ws{}�
�)���}w���Jd���	�t�t�| \@�K4ytçʊʄVrb�4����ߜ�-^,�#m-G#<�1�q�����t-�<�(����
<�$�N2^���/�Ė�o�z&=�Dі��/�4H����O�ݔJbR�[��tx/��zν�O�ے&��M��b�s�.��=<X�A/�,�O�BT�Π'������4�1>�i���-��i��XpĘV0��LA��O�L�N��j�F󜹛	���>��Pۉ�V
���G�pSD�څ����:�"EQ'k�[�C�)b[�bMFi��������7Gc&*JYW���ƀF���Z3.!;���ʔ�Ԟ�\�&۞۟�	'�J(���c8��/A�P�_��*�:M�b�ҡo%���0���F�l��q�i���sv�\��I�\e�6,��AI9�>p��(m�wj����v!
�����z?H�2X�C�9n�������Hl����P�}zk.�{X�r�q������&k0�P��<��Fh �.oU[��L���^e1���7G.��0��Rg��"��%`zUR�K��¹Uh@Y����֢�����$.#J~>�~r�趟 �_��h7f�Xw:T�өΓ|����cW��y�|���G����	TE���p���(4��3�ɘ�p����tq�o����4��w�B�%�Fˤ~���#�g%ד����JD����J�<�#�.�C;�Y�<p��n��i\¤Q�}����z#[M.������2'̼�t�2��CD�
�Chd�D�Gk]��M ��y,°�lޠZ)Pq{��X.	T���wMb�C�6-��7(��O9��7J�j�B�,����p�@���N[�T=��r[i�x����U�U�yiP�g��\���3����
����������M�FC����z���Z�#D�C-e�;$�	�rU?��}�L.Q��-�J��F���D��M.����e�7��A>���)�]�v	P�L�#*<j��Ү{3C/$��74by<)�K����k�4Z�a2���1
�A�_y��	����}��f�� ˿��}ժ�7�a:�ׄ'*B �6�@�����4#��)�^A��� d�p�f�� ��X�������l�� �t�d�k���':.e����|3�!�.B��xpAO=�R�󼴜��}�KJ�M�;��%���V�q��>t�}�m�6��b�؋xp/[2@BV��3���T�1T�)�O�������h�3d�vE�>s���Jvk��X�-�>�][� �]w��>��O�w	81����u	ԅ�A�w�?�Wj�=�6�!��=�툢/�	�(����Y����3v �v��H�1~�,�R?	(o�LF{�p��h��z{��q���ڬ�;�x�����݉X�|�?�3`N��A�ܲ��!>�\��٠����Us^�ȋ�<�1�ё�[J��&D��E\�ܾ�P{��@m���,Q�π4���R��4?^t"�s�z�X���0��E��Į�!4�$�s���}���
u����R�h�ɮ�$�o�;��C�kA���4`��)!����n����w�Wv֮�a #H��� l�����BT/���Z��b��+g��/I��<��Y��D/���Ah�?	8����;�q��\������#�Z7;-}���)r�ܭ���w3'��,.��)�3м)�@Ms#i����Į� ��A8#~X��T9�KcZv~jǴP%�-��!Z,V�r�/z�C�i!�1u=���T�-Q� �����HD[&�Y��9�54����W(��3:;L��@E5�ҳP��R�@<�G4��������ɨ+�664�Z��ÌCD~��3F�b��hT��J�#�µE��s�#-1Y�rB�irY�իs����[����=w��xqdu�2Z� M���V�{�������Z�q�`���(�G��[;�
9�>2¥�E��=�!����q
�|�tT?���GF���(+��!FSAj�>[���0���e�M@�v���[���?A���	���i��\E�ｵ[6y��&j��+6�s���6t�3� 6V�%�%;���_�5ao�{6�x쇦|�w�)����w$��W�Ù�]N�:��1x�.qnDW" N��+�~pt���
����J��Μs�b��c��j�}��N���#R3<-ze�ԅd{Ou���r�dP
���}7j����\?ƾ� |���i�	��x�-~=�S���0�/��}�n�d¸	����A�e|��dE{�9��əY�}g�'��+����=�"��:���6�чӭx4!7i���"͈j����i�p�s�,��疟���.t�g\̏� }#V9RpD\Ky��u#�x>�����\�a��:��(��C��r��Zu�~��2]�Q�Ҿ�FBȆ��h�yE\��ӯ�Ϝ�w�n����JT���[ҕ-F�z7k�J$��a���F9�n7JNd�[౐��t��H3?�^���C8�� m_���nU.᷶����!���H�oF��Z`���K>ں��L���V���H�b��5uXR��3�bH�(5�� �*�)���6����HP�|#078�
���Yx���H�)���dTF��k1P�'l�D�0l׫t^�p�2t֛����O�D"�J9�7��$��[�>���\��˓:��WB�uJ���b*���O�3�6�A��7ع�+�lh�� �I$w%�:��eV�����@ �	r�r���\0��u�!�n�RkT�a��À�1:w3���u��w8@�ٔ��!�=2�
 t��X6&;E��e�������G�� `�t8I�$��ْ�����Srt��[Պ?>[�8�r}��&7ײ�p�U��j�^�{���Nn�� ���H�uy�����{���z �]�;�~<]6��n��>u%�5.P���:�)�v��X�_�l�9��c�ʭ�JxNt���Oi��9�Ru��m����i�2�2%����d�yyב�[v�:Mw�$�r���n��RD�6qi���JI�seT���V]��Y0S�<�F�İD��2g�%u�&����k�M�'�yK�.|B���T�d��7�/|��o)P�u�2 �Ðr���q��1�8�.a)q��%")2�1痠q������ķS��g���a�> ,���i]n�JH'q
����|��	��!�{�x���Mս�U��1Ln�F6��/ƨ$0�(l'���R���Zgg�;ZW��%d}�lJ$�$��t��J=�1���'�.�^F�N~/���W!�>��R�ݹ�(�����&�� n+Yc�.:|�pƟeFta�o{2מ�g�6��>`J���]
���h'���\�D�]�W��e/����ֽ�����;��1ٖ�������`��s:�ּ��_�t0Q�ǳ#(��3���V 	���������7g\i����0�U��p��E��]~3��Ё+��KI��d�W��I_��!ٙ�q���0�<�{�9���t�QL�r[v*�"�daMϯ8�>I��`u���*n��B�}*f��h��%@K2O'd��*���P,�ڞ㑸�7�h���
�wkG�Q�u��U�0|��u�Z�}� �[���3B7Z�ZL��5���^�|;m|�= 'k:��� @=��k^�23
��-x
P����4/^����$�B`�{~�S�Ԥ ��_�UF�b���
)�4�.g��%9`y���%D��� E5�f��~���S�(&#��D��VDT���R�: 9c�[#&��K�S���Z�m�}�q���iYkLy��f3�-�1!p� Σ$��rfW�+��E�.�E�
 \+ P��@fLv��xd`70?2��ڗ9'L!�v(Ƥ�/"�Cp<� .��I�O������^��AW��O]��:(����יx##�-0�BjWPS�$���z�膶���Q��:������u��O��(�ҧEq*�z�4*y�������3:;\~�a3�0]��m�����㣷����ퟔ�h_�fk������Y�T\B��[9Q�Q�'I��^�IQ�|Ƨ4�p�B�lI��	��b�ث��+� �D�Λ|�U�ƼsE;ǐ�E�l;r�z;��E2p��eCKې�'����U
xK��(�_SV׌��j/p~.#A�A�����㻍��*l��R�Nq��K^�I�%�� `*�O�'���6�Sw	w�}�bd:������]j���I�n��õ�p���ĭH?F%p?QX�s��=�Ս�&Pk��� �ilY�P������,MW�.����|�'@J�;���@<���Ȱ���wmrVQq:�K0݉��X�g��c��vK~yh4G+?�j���6�x��U�H�I�~5`W{�Nz���_��M >o]"��f���C���&�/b�&>��	k!�^�RY�]{���2E�������Ɛ���f�هA]E��P�L,�P�@�H�o�:J�Fc��y����N|,~�����3�w�|��ۧT��l�K}����`��M�jH$� PUH�J�ѡ|���'<o������c�>����:/�]�A}G}��6O��d�j�߬�k��V��Wؐ�8��u1��a�j�z���(:c;�:�s!����Oث��3x�>m�J^���e���AB�9�Z�R�<�/҇�[Lo�V���=Ԋi�H�4�]�T"G��n�L�v|,�Y+������1)���U-)q>L�/��A� ���gH7���YJ7���O��7�R�f�w撷/ؑz8��ē����~�z�e�@ik�����\�.���Z杆�*��:��bڟ��������
�U� н8���@�.�s�g���;�L���RZ$��`A]�E<�T����"�Y^2�d!����[�~��m�̅�s��L��"�A�%�~Ѵtf��E���O�]�x���>�pjd|<s�Z�z�W�%ԗ.� �cZ�i�9	Y�d5��9�W�u+�� �B5CY�,v
�*5��J�4`�9� e�����.ɑf��s����B@N1� �%|d��vw"X	Yj�ŝ���*yX ��$.f0�aA�	G�Q��7>��Ca����S�l���j����!tq���~4��k��u}�>��Q������߇�����Q��$��Ŷ���|)]m�2�,��|�̥$��g0�l1@�6ڭR2K�.�d�s��QhW���Y?֤_<�s������1!�wG��	��h����POD{�ë���vbn�j�4��j������|qWG�R�<Ҩ��g�ƙ�Vչ�F�?)�&ALfi�v��j�~��W+nr�-$<���Ѧ����z�Z\(�~`c77'�ⵑO�Kܕ!���n�EYO,���rP�?�]���Z����H�9,�B�*�p.݌��u[C�yʠ�^Z+?��$�;���z�9rl�_<e�?ū(Fo��!��%}�rg���yv�f���Uf�����ͼ7cϹ�F�|��r��
�S$#��p�O��I!L�ISp��Jl���pX^�17�&Z ��xv:�T� <6A|v���>�b����{i��c!�$����Q�UŝՌ�{� ~�7�)zcХ�65<2�����F��oK5T�&9�C�XM���z}��n�g3U�\6'*�b�&>��.[^~��p��[��~�@6���L�x���.�â�W�[�#�/h������Y��m�5L��k�ӏ���2!a�#7oM�Zx�%v��3b��q⯐�w\A�ͱ��T���)˦���/�2D�� �hpz��t� ��8駀E���M�/ =N�y�K$�|�l�(HF�U��xn1��������'ubN�c��ge��T��C�[PWk^e�hy��s�܄yf4