��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]rܕ�u���4�Vrnn�?M��Ov�&���rd�\
���)�+�Q�&�����3-݈��Vq~��MȆ�W�����zŔ�+�n��OZ���vf*���@Uf�M�+!uH�M;�*P���^
V��#K��ΫW��:�N;֚m'�a�jJy��)!�ޥL7�����ˠ���%����=���TY��̨aO3�[�=<_XP���-��Hi��2[�E��N�"E����C+*^kҿ(�t !Z�F֧��3ʞTw��&��ʧx��RNj���OX{w�M����	���P���y��ʕ��w���}�������zL3y���Q�O�բ�aB2�C�c�=�u��t�-f�%\����Z$����K<����R�~������YvX�꽧1��p4���5���F��F�<C���~v������2�k��a+n�W��@ֲ��X�wFg=��L�`�qsb���R�ǳ�;��g�֋��h�,:��j}���}F絩W���n��$��zV}�N*�A�wJ*.s�	?E}�`%���l�Ƀ=�
�
!��%�!IV��^���}<2�PE���:�Y}	pL[�Bo0�E$Xn�(�YK��.@�R�ulό
�
��b�H��PCx��c�:i��߭G�[Zl���<��9� ��K;��yMI���s��{�`����[L�5UI�٠uф�c�+M���?Q�����'�U8xM4$���v�~8'TJ�M:�bg�4���]<�u{,x2,�趀�%�B�O	�D�Q���C���B$B�Hs�)�*��һ���.08xk/����r��<�LC)�	��7��%^���9�Ke�-�:W�S��}�\��D3�hA)����9�S`��ѵ�>F �	�Fk��+�
��)w������e��Ӫ�Y��Ht�W(I���PU��u��C�gȨ�I�����~��9�81���v��yN`=��+��V�Ϭ�HQP �
���֋�(�����n��T8� �"'Ғ��E����m���B��b+����i\�c�*}�"�jrQWa�ױ;a��tamzf`�{�^�튰I8�)E��­���#�K��5�@��~����u���+�{�7Q��&�k�����8�B���N�N������FX���@��r��R,1��%�;��G!`Q�ŧqJW9^�h�:���-U+�j���Z�p��,����Nu�fϸE<����I(y��֐g��l�Ev�Q{#(L�V(�:X3�Rw?���*����~j�K����`-�����vm	�PY�q�_^�~;���4 ��p.,�z����Sŵ�=��%�~J1��\KU�Ў<�Jq�/~�j[����\L�=4�ʉ�M�2�0o�sε��� a�ۆ��ߧ�C"��%���|�	2`��4.�30��;zR
��S���l�Ev���^ˍ�6f���ѩ�EY�:�2�3��W��j�ȕ�=�cY\�6�����6C����w#(8��Y���X{o��ID�t�wk_�}�W�kc5#R���ϐ��h�jF\�����o���n\&v���/bk{r˨�*#�*	U~�>Y�Q_Pt R�CO�|;] ��Ov�W���I}�X���\j5It�j��|�r�٬0�eB!�zm�F���qX��h���v�7��KR��2%GÓE�X�+Q�y'H ��&�%�m���ǽ^:�3��F���OV ]�y��ֱ��a���Nm��}��^u��0�����$ex��8/0�hV����_h�<N�3HT���P���%�r_�T��|�&��
�#�IEȺb:�/�Z�,����
̣߬�<�o��m)~ȯ��HY'ȋ)+84�������4�+cǦ��pe���,�Z�1�Hm�����B� �MZm�9��7\v��ʋV���.�]v�Y�a��3e��W�?��j�DK�c�Þ��̘�*�;%l������<i��H ,��>j$�N/!�n���)��u���-X)2�_���6��j�uh6/4*5�
@, �B9}7���I��U}8����N	��*-�#�Z_!�U? ��JP�t��(+]j�_�d�Y�����u9G/2>���w�o��#T.	��L��}�x΄�� �j�F�1��^�Tn�g��Q�A盶��.�.R�nme�M<:�F���G��($�v9W�ld�7=OM�-!��J�����U��k$��T�8|�5�H��v���hQ�-/���?�m�k����:�$P�];�n8t��T��������&�j���-���+�|�DVd��p O��6���RS'�e���e�Ep���$b���+�K�{4��pq{�e�����N+v8�Ƞ.F�Hm�!�k�DE#�����͢.p(�5�~��.�`,���,��g�[�AP��<2�򽟵��@ܽ�m����摔�����0y4YJ@�:�ج/6$c>>�0�*�(=L�Ǣ(�-).�%'d��mY`?')��ֿ�����s�ո�ET�1aC;]>���*E��}m�à�x�x��[C��%��T�_eS�B�8�HjUpM�����j�N%,�F�� ST{���dԀjq��2}�ūD([�g2�4�9��Nf�Z�B$����f�[���si��E��Ӄ�|#)��ZrPy�����ݽ�>��5m*�M�E˖�2՗�{�9?oBD��Uk�c�����̾�\�e]*����6�H����Uϐ��F_]�j�?�Xf�����ɐ���	�&m�$v(LE��&���z������@ݓS#<(�d,�D0��R	�iΟ" �P�$z��Q߀�2b'M�,U�`Ej��5�;D�[a
��;C̴�r?�4.�o�����%���gPc*�����+���f���D�l1Hi�S(J�C]%��9�9�3�(���U�0�4ۋXx7�XMm�t���9j��t�1�
UD�N'u'�z�u9b-��)uy��7c�͝�ե6L��J?.z�Ld/�90G�<x�b^ы�Z�)O$��c�ؙ_*�Xf6* �KV��\��r��m,>Z+�#�m%�e���\�Z��$��LX�:p}Tg�I�����?4	�2Sxy��a��ecךs7��11���tHC?FRJU[�Ay�����ѷ�B���+���7��X�'z6LF�qG-��dV�1�r�݉�%�Oj��,k���\KG�0ZHm�^��}�#����wCS�ěo#��&����+[4��?�z�*;��.�<�-���F��*�0B�`V�;�H��w�0��o4d�'�-��,g)=��Eu7>\z�緍۩����@�|(�%�����\f˴ҕ��G��Gީ���&\���J�n�l���a?���f{\=��y��V��j�+긽�d�xL0��,�my�$*܀-���.�1S��XGR� ~[a��ܶ���.k����d6��:K`�|�Q��
`OB}�l��Z4�ŻqL~��?�F�F,�J�Ke�X�o�2�?��/,(-�'�b�&Hj4D��<���
z6:]oح#�1����6(�Q�$�� �p�~?>C�gϦ�ʃ��d� =q���g-h�,��Ǌ]+FF�U٠Ə�;k�#�%;�pŇE@4S�n(5��ȓ>�H��F�I}������;E�����#7&ER�4w3GE��Nd([+g�&��l�W��?�N+w�:Q��^9�����/�
6[��U�|����B����r���~7z����o�I齆RxH�tn�ʍ:���,�J5%v��@g�[m:��_^�KuƼU��Q��g�S�ZN��!Gۊ�Z_ �~��-u��8�3�����ф��N�S�_�<�M�D��Z��F�l�m��X�.�����`��=�CY�jѾ�M.A1/���O�n0��͛��ʈ<�Ҏ�������yz�G��^/[������8jR+ Ic���P]\�z���8c,D�s�t���V�zH�&�8~kFl�"�c~S���=i��Ԟ�<	s�ߵCҀKT(/�d���d��0�p�p�-2a�m��)#Dn.����ѿe|����&]UN��o5eE����L���ʆ������
�����jV_�7�G�S(u�M;�ʒd�Ɛ����|I`Z���m|�&�Zd#"��B���k��P�h Hf7��L7Ю���٬��͔��n� �c;�|ݬf7��Hފ�t���d���WL-��5�D�i4�j*��	`�Z�����r+�Fz�Ayiy+��'��q�fHWIӳ4g+�s�gZ�}�F+&�3�d~�ɹ�g W كN��ȍ؄��-|���j[,��"�KN���sgN���F%�3�̅����dYW�����us���⤓��s&i�yh8��&�B-���Y��R�?���ޣ�M�����:�Msn��%��%6*����)�㑮}�L�X�E�;�����>�b	�������&_,q3���?U���{�f��/뮺�~U���1jv��+��޶�.����*}�Ov�l�fu垦��{�xI��=	�en`{9�C��~��!OЪ�$w�|l��.Fv↟��^����U��A��}pi�xz�r��������g�i�$� �ƭ���es��V��<
�GiJ�+q�7��Lc��m�	K�E����Fj~\V,$��9�I��C|͠d�n���B����p�[�sf�@���IR5U�g��ѯV��|�"6�3����b�K��U�H�u8�(�oZכ���*2x#�dXN`9tx`����W��l��s���a��+[�[��x�B=�1>��<纟�}�-�h�<+�^���1������b��$ 
�@���m&gci[�B@1��W�ӆs)wi�#�����4��̑���a+����(
��`�6�]���x[��]��J��j-�oD���z~hN����HQ�NRe�{۠aS���K��kĭ�$�7�O��v.�t���#��[��cO��~�Mk�dݮ���y�����ʷ�-��Jā'�f��h�0�ٝ��dgU
ˉI��deQ.�8@ӐէE1/H)��<�Г�[�'�M�g;nH0J˒��r�-,��òL��M�8�$�o����,ri�r��)D��o���֕�s�X��v�/�%��O>�師�i��z�[WNe�?�`N�u��5:�1�8�VY����&:��iu�Q��_%L*�;l�Β�P�٘-sݵ��?���'�3>���tX���s�i���6>��Sz/<XFϾ�n���`��܏��� F�d�,~���{�X5�]r0Ǒ�1[�F5���wwr�/4��y)���'`6��>-#��KJ������H�W��ԾT٦�k�ϻ�ך1��oo%�:�ZxcqY:�MN�Nh	��	�� $G��k7n�?�*��y�\���7����]�����\���M�� �13���Y�@�Q�"w��V�zͳ��6���ӀI9��=���J����E�wA�������S_9g�����f`4�/[˥�:����Rqp��
{�
2�'}\ά�ѿWk�cu�̱`�<d�$����e4-#�!I��w1;PO��k��Fϴz��s�z/n�ms�Ǥf�c��l"*��u�7x|��c[�o`c���T_��@�R��b�ٛe�,��u��!hf|c�0�Q����1 �;=>F�}��gE���Ƹa�����}I�u�TO����k��R�2S�#�������|�B�Sm�(���t۲���T(�������;��B�c�J[�Ц#��M��u��Z��G�� �fh0z$<K0Ni
A��"�K3���L�P���S��p�H؉d�A��F�������r��hMo
C  c�t	>^�ɨ���:�'�\�O\`ѓM.��e�����x�����.���)�F���N4f�_��T�����gxCq�F�̣MmT���E�"��1I5e�Zk5�2�u@�����A��8p�������ƥ�(�5dp�r��0WVa����Yv����'���ƺ}[q��"csM䭯�7�b����Jcˆ��>���iR������3���9���hWh������P�?+/$��L�_L�"��i)f^{�@[{L����:�[�W/��3k%a���A�͂��p�4�����	��0�R�c�~�Z�+&�Np�������T*F�܄gp:�eR�ʘ�a�zi�~?t�5�*t��r�a�$/����݃u}��wi�J҉��o66#v7�#B����߈��Dt�a�Î��lf�d�o��5��d*	"�����M�W�BD��2z�x�2 ���-NCs����W�����D8㜱�7���V2S,���刃�~��]��(3 e��!�)��V��3��W��$�Q�u@v�].Z�$6c}�'����!sa��^0,iPzv=��b�B�X��j��S[=mz�_;"e�S-�kcZ��(c�U�I����4�S3� �@{_�䁽}�VW�;�S%&:��/EC�H�����<��&ц�� ��sZ��_�*@N�>;sT�b��Yδ�x�dp�X�?K�Y8����
l�P8�~���a"�����1�PK�(hб���+Y�*�(��W��`+�0ع%�y4�x��g�:O�����H�t��_ �����Z,��-�!����Fyf��t�@8�$n���^'�Ȼ�"���m[�ϩ�~����Qn���p�����	vZ������<��ͷA���^�'�(ߜ`T��O�*�~AeA�[2�G=Z:^~�Y��FT&�Y��s	 �$Ǝ*� &����56F����s��MNyi�t���ڲ���ǫX>#:�����W�N��߶�ut�+��pz>c�,+G�/�zS$=o=Th!��lo�]kB@�����ś_%�C�>'����E�6_��e�����?�U�U&җp��G������Sߔ�����q/I� k��vF�DX���Q�����`��h�q< e�a)�&�b����[m���4�Z���~��:v�2r�{�<�����U.��o�6f�1�3Gj�FvO��͕r5t�+�'���޼�!c�NR��~�Y������ܫi <y����jy�HBqb�KR��;���8����ٱ���PQ"|��9�V|� ���=I响�y�G95O'���WN�D"�o�;�č�_ƥP<�IJ�J�MX�8:S�!;}�2��K�Ņ�ב�ݝ�Yܯ�	2�|��k�o>%�G6�$�ݨZZ�/�$��0Q(X�������P;�~�=�]�z��QU0gGL= W�Ab,Ӳ*HO7�($�Z7g�������7�MB�ШpZeC���Yڃ���'
��p�����x*��@�-x�|�ʐpBGecH'����L�i�=X�\s�Pub���d~l_��fqj�� �v(��d�^����I�z�^��P6GZf�I����Y�+��\�ö�M.'�M!��>������C��i"oT���X���l��*e�@�1���zWh|��D�&߃j\�l�)�?s��������B,�U>�ْ�!�*�W�v�۽�%��q�{`C���xOS�b16��L�4|��ɧ�dC�Ñ�>v+�ͯ�g@��M���	pp��p:;��u�9�䢂�Ɣd{�Fùx�O|��!�Ξ�[d��I�8��%U��r8S�GÎ��p�D{[�"�װ�d�H�a�����R��ڱ����:��T�p�����H�f��w<P5�fn��޿�]rkop�"9 ����O��W��r	1�ɔ���Ż�����0��D3�i�"y�<w[9�����p-�e���~�_ �)4�4z�����&+��i@������G�ѓ�z�d/3�����"��C�4��@�#w��E��gʺ��O͗�(���e\���U4؍N"���"J��_�p�[@5&�����s�(�S'!��˯N,�6-�g�]���Y���cIf
�ȸ��p�;��qu�R�Ի9߱{��|m�p|�D:���L���0i���l7�	��N�=�b�Qc��8����z7�tbH����JP���Ռ����L��K���|�T1bm���8��N�nN%7���y�8��k	<�Δ�;dn�B�0���;�v5e�S0�'� �0#�I).NԄ�,��1�Bq����ĳCt�Z]����Ѿ��C�K�W�����>��R��6b��~e�`z��_�(C9e~�8p�3��p_�C����l6��O��C���-�~�!�C�mI]��)�U�[;~Жڲ�,�O�������"d�?�>w���j���L+!��6P0�mH-y��9��9i ��*��.
��*�� <9HZV�
	�����Ip��Uɀ�DDXU�"��X�*4���v�{:T���<ƙ��ծ�4��v1�4S9�Oy��T'����Y� <�[���Ǐf� M�i��CDk+�{��	�I$'��D�F6����We>����,h6�JӁ���D���3P�rUs�mp�SC��I]V��M�mDy��y�B��ҹ�(����k��`�4)�\�'�` 0��'�nLg���?���ڊw=$��r�+�" +�ٗt�Ķ$Y��Rv���D[��U�,�q!��&Ӏ���36�l�*j��(7 �ޚ)��M�?��
�r�� x�X̵>��:��D�n�Ȩt++t�i�z�*��x�\5�ǳ��O�Ip՜����v�z>��6:՗`�	�($��/ִ:Ax
��@�!,F�
F��2!Z��:UA��/�?ŇO�������a�~$kq�v�	j?�iUp�Y����o�j��Ð���	h�t��_���o�U<���u��h��@]��CZ�ןe��۵	�Z̨��c�֣o��Q����u�3z5�n]������<XVh�C/�����JՑ[�p������Y�X�+P���F����̐��O�Ĳt��-��SC�O���H��k�|X��6����8�
G9�(*��cH޻-]��C��p�u�v,�$*�:��Mb�ڠ֛�p5OXR�(05�ӹ!��SC^?�(,N�@��t��"�Ш�O�v\P��֋]�N7'�C�쏢�Xa�<��;CdY\���ҥ�%�qʼq�;��b�F#``�MU��+��Y��,�v�:L���[�-}^3�gc�����Oh 2k�3HT�sn�:��b82�������,zJ��4���K����B�J!w��G�5⚵��/[�*��}�*\���˩P��.E]����vg�u��x��z�N`�t�lyv���\���4b����*	R��H�W �ø�s]�(j�c�V�Q�B	�.G�&�������������R��F�5�AJ�o�Y�Q����Θ��o(h��`���"h(�Bd��T�l�Al���-=�	�)q�8�kHظO�ܴOķ����x�弇MH��R��:�R��6���[0ݟ�I�(�%-���c1Q�8�C�M�������G.N�dT�]���g��~%���c�-�����D�݃O"6aM�_3㨄�/�]��[)D8=G����ޤ�k�1��cYl@H.��dMV������F���O;���z��3X�; Q[g�}p���cQ�]Zg�-��u��q�H������m���_G�{�i���S�u%j�G���i/��?+��|�[gd���0#ǕzrD�e#F� /I�`]G�����\�O!���&�U�� �ON�:cHg+U���5�e�Qk�/�_i0�F�(����#VGmV �Y�#R�&L���ֻ��L���QQ��ݪ����N	D�d�5�~w�5��TB/��t�V����6Ύ��I�Ȟ����-W��]2
��!Qp�Lt����˥���4�15H{SA�8?�>�]��A����A��<��b��s�����N<_C� 5�=�Dd`8�ᜯ�۝��:Uh�I�M~C����*h�-���7�m�C�i�</b�f1	K�d&��|*�	0�gx��4��!D�ޅ�`��z��>bv�H�	0/X����e�T�~7�n�٥�Mj_��!!���c Fk2&h�Y�,�3[��_�v�g
����;�g�3�Zb�^�
n�$�`���<�)pdı���O����zX���$��ư�@�@��k]G^LfB�
��D��ws��0S�%Xҙ��#����e�(���'D�-ķ6��$ҡ�M�qYO�I.�!n&�o<֢L�(������8�n�TR���kQWw&�*4��[�����}.�q���G��{������a���0zv~������������I���/� Zh�[��x�C�ڲ�)=�,5�ͫ���P�Q?t�P>��G{�p��K��2��1�)(֝��IC�B�I8Z�!���+׻_��{bc��z���o���q�L��ctW��a4+����JW�tI�a��hJ[�|�Ýq�N�j:c)��i2��@`�˥�P'�:	�ҕ�Y�m��=��FΑ��֑��?�� ��/}p�<�<B��g,s�R>	@�,������Z�Z�j���83��"���pV&s�ܥnGY����� vƟ;U�
5¬�#yZڤ��>V��):��@��G�"��NX��Z���i}|K�!�s�=ɧ1L����	�G�G�_�CBn���B6��Hm��xI5>nΒYT�S�Qj#m�o�_�_aW�������K�w"�go�H&:e@M?��fƲ�gGVGW��e���u��ym�(�,�ڿ��t��SX�����.��G߯���8�Z��=y�V��>�4�˾� ��7��S<+3L����p4te�����v93�P�v�"����Y0��	p=������M-���z?t�T79�a(�!�K�z�	�6XN��z�g'��+�{;�]B���#V�W�tԽ�Юs�п���f��S_!�.~���e���[�[$���\J�ߌ���
5v?�?^&$xRM�K0A�0���x���{\0�B���;�+���lٷjzN�@+�=��� �����Rvi\y�����W9��i_UV�6��?�X,0��|�z�'�5�a���卑��tc�2g;�#dI~��?���~�&��'����GM�c4�Ӏ6S�ҜS��6�Y_������Jq��J5T�\eoB���|����r�bZ�4��ӂݴ$=�������� 9f��M�T�KYd���&j�r�/uL6ۻ��Gp��TH��BR`���	�����C���G�B[�t�+��ޚ�48�i����h$H�oI^O���u$s��'_D/�LC;��]���<�L��g�Y�"ã����=S��ʚ�"��U����D�ߓ"��}�2'y[(��R�7���p��^#8��־��i�,�. .(վ/(����$�{�ڽ5�j]�8�4��զghPCњ�g^����7��wz4<�v~)kkA���02񧟟3�w����0�����A�7�C=��|6����(P`v��Ml�lj��s��r5#=�ĭ*"�����D�bew5`W��Jm��ͭ�bؾ?���&�޺~Z"��:��O�@���Y`�� '���&��h�������q���p�NM�M��/I�pQ��'���6���d6Ч<�P�Pc�QF]��s
�P���nн !��j�S�a}8P�H�.ce� Ϯ���i"BǬlg^�ֈ��p�AjO����	�*)�GgqLp�]�-]�Uku�`�*�"�6�&���n�^���f�˕�����f�ir~�f?�n�&�S�>�@n��|p:-�]����]��t5۽Q���U)��»Q<C������5���R׬���q�r	���j�wL��Wn!"����w+��x��)'E���R(g3{k��qN%�+��
���?�%s;�<��� @V��o���Xƴ�Z�s ya�!�1���J>K5��f��M��HB/']��r���T�`>�?4$�CO���?@�
n���=�o�`W���(�S���7i�Y�)l(^�$ ��p�J��I�G����z/���)��"BqZ�-"W��x��<�Hҫ\��s������"�V�'E�yzT����q2>e6>z �Á�ݝ�¤�k3	ƼOǙ�9�~F����Q��(�s��oE�L�G-��)@�̽$C���r���
\�_�nݒ����OzcO��EJ�<<��2���c
�{�يd���%PK�wD���`8�cu��2
�V�����Y��n|w�T��!�Fc���p.���~fw}���ډ������*L��Y�b,?�����0���7�J�*RL�H^!�HJk���n��gR�m{��~Gq�D���=���`>ّJI.C��c�Wv��4ä� C@ݑ3s-��\U|�H��<�;%XI�m�2���f:��#��l��l��E:���e��8)w�5;�B"���5ݰ�.z�lr�:_,��R�s�$V�����q�Zh��f�*�H��^(K��p���1���d�f
*~*ٝ��z�����n�U Bw_1b���QN�K�B��RZW��2�͠R7ޕ����ן`�u}Q�i�SI����On:�����h��
"�	f��k��=d�c����[���]�ʅ��Cm���%�I_0z�� ��sR���zy�H�W��$s�����C ��v�q�{�w6�rW��exCW�%26&IH݄