��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su�XT|H����y�M�a��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P����3�T'N%w��d!Q1%�7̬�ONMς+���u�'" ��)�4�.��R��L�0*��vX���Y��EY�U�R ة`����Iʘ{�Y*�b>����4�*}y�:$��i��-7��C�I�QPdN���� m��3��=K!�3 2��H�l�8F|��w����5�i؎���"�^�EX���m!�W����Z�:��:�=8%��@���h"P+������J��<d��	���J~�-��I���l�5{����Wa�W���T���w�})G�2H�p��z;��-��D|���z83�8�,�
^N;vISt��.���MOl�c%����ƎT�$8�JLGS�(T*2�xy�4�2��]ႎe���ۡMǣCҸ�\z���q͹4;������1@2��z̅qg�~�ǇY�B]��g|������cۑR��4����oi��_�a[���)Vp�g���=q�'��T����g�y�=���Z{���k��!Һb�?�~3��5Q0�u��ɞ��m\�/��U,���Q+'YJ�,���D]�3�H�~��@C<o(�)K�&��A�ֿxM}� �F�zt	S>欄��9�%ڃ����GH;h��P	��2p�yo�R�� �9�E�,*~���l�1�-9�L�c>���H>�e-5��[ot2�� e�P�����A�y/^I�?�}S�:�Y
�~⊼�?����y��i��{���ʽ���-hJCC�R�6�}Le���G�R��
X;�t7u�>HڹV��2'�o=�,�'Zə9^$i�����&�������,/���Ь�R"k�9� �{ޟ��� ��D�\�]2@#F�������@��r2�3p�x�x��l�	Z����ܮn�W�.
�����Ӎ�xX���J#	b��>b�t"[�o�'h#���y�!d���y"�w�	ț}��#��S����^ɶ�.���5�u�iY�M�(w:#]���꜌nU�'�V���<��>�%�L)b�3����-y5g(�h7!|���v���b�n��6)�U��u��pe�xX�c��gi�痚
Eεwi���=�K9�ܝ"�#${��m;��MV�Ōc��������|�E@1пԄ�����L
�_��i�< �>nFe���eQ�~�U<��Ce2|!��!�K�"3�O����T�I�to�������a��������.��6��T��r���4�Uw�@��S��<����e���E��|a�m�P�t�y���s��8�4�D1�g�e�p�ham�g��@(:���u��13���EŨ?���ѥ�P����ˀ{P�g�Ȫ��Lf��V�W�J�"�>刴*Q�ۚAt����2\GV�����	��y�6e,	��_��G�Fu쒭`d�D�V����q���Q�G0`7ȋT��̜,i��,��I�7IW������7�p��2�zu��ˬU��b#�=Eבb����[IC���< y_�F���<�}�ѓ�z Q�CCT�G����bO�$`���/��%�j� V�6�| H��-D|��U���#��X"n�l�^�G�� ��H5��Ͼ]���8j��g>|�IO���{��3�D�K��A��w>�=ğxh���������e��x�"�K����)�'�b��!n�(���y�5�P���B�T�
 8?�́%l��z��xv�~&d^��au�����;;�uos��剿@������H�-b��QbmBX�-F}5�DF��٬���Y]D��/.�	 ?9�t}���]Åg-MBRa[�0�V��	�s�u]^qq
�4[�ϒgu�/%o���c$����_�I�7X�����;1��?�K9K�hF�����:F���gP���U~?g-	�)����N3�)0�@�L�?p���fHv8J���cȭ���< ��1������8�ͻ�Hx�/��_B��H璼�C��e�ɷv���8���.h/�&�!#�K/�����t�|	@�67)(O�ȵ5����*��C��y�5u(�$�A�<D_�ճ^��N��a����LJ6���w���ѣ�5���sz�f5.���Y=�{��c�H���M됧�tH���"���l���}!�#�R��g@*r6AL�;�"��H^X��2��Mʳ���ԅگO��B� �:ئ��a�e��zuRK�ew�Z�x�#���� �ԭgOC��A�@ XC���|ok�D� �R�h
��7��s	{;��01M�|?x��uyIm��,��`���;;a������z hf��ˮ"?�(�z�����ה`�>@z5k܊xD�{�қ=�fޤM}!~u����C2�C5�/� �ګ:Ħ刺sY� 
V�	��!��!a���A�8�|y�-<�s@�X&}����7�f��]�@K�@�b^�m���K6;��@�b���;:]�7�W2�v��/�s"E�}�E����B�4"�> �Z�)v��8v����k���حpz�O�W9?y���R�.α�9��^l��&�䜾����Y����?�njr_j�2 �]n�9������b���7'�+8�P���X�҅
���51#G�fT0�%~��X�,P�6 �A��ׄ2c���\3�D���a��� �93�	�G����-�{J�� � �����􋀯	�%�Gn�tyi�C�c���s0Ys~�j8��CO�jf-�y.�|-�r��Ko@��ɟ^~�{�[��M�7����$%�Z��t��P��u�
�0��!��i�
s�l����+���DS�C%�.�ؘ؉eB��%�	���B��.0�����*���|N[;2�#���_D�c����n�օ1L�}�e���=�[����J����-%��@��|�Fɜ~�*%
���%��`Q�1~���?9q<~z��).�Uh3��>֨VT��HO�ZEYk<�
�B���`�TuB�|:I˿�{�beb��<�#@f�2b\j|<[�BfB�H��&S�u\�]yzg���\z�$�(f�Z�q��_/bd�~�%���kp��	r���i��p!��2��H��tI��φ�������B�����dJ2��V��Μ*g�['�s>@��W�V�/ ��A�/d�9��&�Ih���kj���>/Q����qy]�s�4^-�MJE�*��Ң4UmͿß�ˬQ_ֈ��*�(.��<����<�7kb�|̍=}�}�n8���!��E�Q�rnvE��p�G��|�3�ezLX�K����>��s6=�����y�үQD=9ã/ŷZ�j3x��o��f��+p��c�a��
q��a�Q���v\��-�ӨR(� �Q�z��d겷r������_s���[.Na0t0�b4�I���� �U�u�axG�%�)%��-��c��Z�_�0��7�6���vw�H~Y�(��VEC߲�*��ο��]k�갦@@��>h2!�:�[ZM��kG[T�?Ҧ]+��k��e#�^� .�J�;JKQA��3ׄخ����tV�CJ�B�И�(��Q���T��SM�,�;����,�80�1=R�&7��6wA��ʮ�\=�w���oEؔҟ�Z���t�'�k�a����ǐ��p�>�yW��M:��j��G���!		B�F�/SȎ�x(�.>�g|�-z��X���3q��j9��/v6 �
1Gb�
Xr�ռ<��T��0~>Kv�@�gm�awg�����[c� -�1@��b��u���DkR�V�&�+|!�pc�*�u=r?ǽ�?��d�c,}s�T��A׃H�zX�E��r b���8T�,��અ�h�~=����4<o�;��Y,�e�3��:��V��Ò%�,���,1ۉM=���H�Sw+w������_�� ��F������[m���WװA�K.�O��m�\�g�7��<�Fyl���>�%*��|v�*o;э��d���c��&r�@�XΑ���}�7�+�Р*$5�>���o�gV^y,޵+1e'],���)+��K��l(�C�+:Nl�b����l2�Y"k�23d���yݗA�q��c��9Z�B @pV�S��!��;xf�@@�I
�G���E�i���Qԧ�$m^+��FV�����<���L�� ��M�إ���d~y&<3]�����UH�P<:�/rjg��ƃ�����=5��G(�?��N��G7��/���<������ǒ��F���!�Ss���}A֙���K��JZ�1�C1b>���l�Q\9+C�1�?.
�g�"����M� �)e)�' Y^j t��A���cj�Nh�Z����"(f�O�{�ʷ�L{�R~z8��U�.g���y�pM����^s�M#m�PM~�j,߀B1��V��,�*f�=��˪��R{���R �V,|�Q((�埬YO#���5?nx�=�N � \ў-:UHLZy��W��[�?�� �s�(�����~è�q�S)M����g�0��?��C�����z.���y(���l��C�B����/���Y(�q+�oz`� ���w7�L$���K����̦�sJA��n�y���y��(�aYδ��v�m�4Y[qK�Sao��㣘�R��� ��	�/Tc�b!���ĭ^���z�m�X�O�贑���&cr�}�>]J}T=W�u�xt�B������\�-d;�q�ـ�N����F7Xk��hi�	�PgZ��C?�?�Z O*��������G8�~nL#�zV��ж�P��
���f�m����/B�}��n������[J�{]��駒�[�W�a6�!Q��5�8эP�j#]�3M�ݶ$Қ�1�$$��rq�/����j�p�`昅(�ŗTF��p̏����.���֋����]�#�8S�P�Z�\��Z�'����h;�<w�0g����0��t�ԦW[�����9j�����E�LR+���}��аE�]��gTE@Rc�{ns�Y�j���[�b���h���S9��"� 뼛!�KH�,|[*y��1na�.(|6ؕ�\�4���L�[���E����9���,J��ީUn2c?SŐ*t�q��h��.Ьz�+�+���҃&ɔ��O���O���^_���H��?��HW���N,��ݖ�9���`�y���z�� z�P��u��:?:V�pS4�˵8A��N�.�'�����5���2�]]@
���*�X�f�������t��:�أw��.�(��̴�?�F�u������ѷ�6l�3�Ύ���&q�M�Kr'������;�X��uXm�MOS��,�z��š�Ps�on�Fu�n���w$�'��qy����V��.�[�:FQ�x6f=|����!kAS7i�0?������v{�.���Z珷�K���"�$��.}<�:���^�2�� ]j�z���R���_��Nw����AS25		t�%+4<e�Tk��z��MU6nx�It��|̓�z���|��x��f�z���:C�O!ޤdXz)�ֽ�Ya�4���>�ģH��y��&jhP� �U�N��ه3��9N9"���`�E$�<��)"0ia;�8�Tդ%�3�M嶥]��yx�i��g�2~���X�j�~�z""vZ�>��Sm2F;�t��-�~AN?6au}���d�� �7�B�u�!��+�_wZv�֢TD��d}�5~i�gWcT@h�W�b����A��35a	�!�f�uBl\��A�9T j�������P��K���O;�W�K|9+;�_��bt'o!q�%;⎼4��X�%-GEs; dY���VP�Mn_�s�����)�!Xfz��E��ξs'���k6i!���b8g�]���C�����{�l"s��C�n�CμK����=����"���}�	th;��[�X����ZQ"Y)�����y!W�fa:n=�P�t���4̘��e�~���ʮS�7Z�ϳ�C�i���`d���(��6�t�,�*ne7���N(Q�����E��.�F�x���ʥ����3Z!%�u���nl��D���x�U�z'����DH�4ѻ�+��D����䈛j&��	���;��b�ݺz����S�M�*�y���J�#Պ��w���Կ0Nb�����A)@�,5fY����K.��K�t�$<Ұ�*}B���@�&F�Ngb2[.�#�
���|�ꈥO,l�[r���<�K1�H� q�<`����gH���a�}h5��D �0��(!S���m���幪Oԫ�|G�#%3L�fE2����%�d <#sB\�s�6G�G"�u�|��Y���S$=W+j]����{��?�}��3�>�L+�`}�ct�N_g���WI�1H��Grbo�RSf^J5K}϶�y�G�K�Z]c�rD�6�)��h��=�@�4LQ�T{�N8>��f#�h�6�[��5C�qHN�uM��R[p/H�g�O�@z�e�Ŷq�(��E�˞���~�M����2���e�A����a^��.Y�ߚ�ح#���{2x\�p�8O����-K(ۍ�'KE�ZT��*<�Tp�׸��n�B�N��"���4M�*���}��zfIdO������Zَ�e�UɻP�9K���p��m`����l �~�:�&����.�1S�4H��W)�do�쾁�(_�l��)���5f���uf�*%d��W�k����69���0��Eu3�8���-6��a�߷1��G7z����(��
?�����64*�x�`'�aI��t*���`3_t�����7'x�j֮�g�.TBt�>��+�"<K�6nw�ݡ�����R뺋�~�s���;:$�G(7N�_������vR���w��`O�}��p0*S!�v��Yz�xj����t�K��k9E�]`�G 2P]�F��n�lݾ�Ҝ.6��)km�,<ӯ�S�~a9x`��7%9�����[�M]�?��Y�Pf�5�3�T	�W��*�~T�w)�@�1�9�E򢰐j�w�%�y���u	�5�rY]��>�n��ŭ%���jƙC3���>�xnN[�����_�/��K�sn��!�g%p8���F��Tg��QH����l(��)v��(�.�|�]�i%����W�`&���oڢ���� ��S��C�@�[�D֫�M���C�����)�[��؊�9N�lT`�4�_��[wym?�%��+:,)�݂�Cp3o����%�_�x�G��O��+�����R�u��V�N��DQ��l��/Pe�rK�v=����-$+�&�x��%_(Bb"i�])@�;�`!�kM�LӃ���&�"=�!���(=}b@����V;hMƤ�x�[*���G�6�5\c�mmx/l:b�7���g����3�;��:� �����CK֣���8$��}��+���ǅ���Oa�~8���Ha'���L��&�h��N�D��ī��PO�,��Hc�?�-����fb�k�AyLfUi�������� �9�]%��V�,��,����w�Ջ")��D5�\�������9����I�Kq%�
>D�.8Y�߶4��k�Rc�U���'�' n�|>��n�P���~p64^Km�m`!Ph�hvz��Jo砼��7+�CŎou������"�l{>q��a�b1S�
p��J�ߠ����ڏ��Lܖ�w�֌}��>�[��
�K��"��9t~8e�l� w��:�Q����dѭ��]�%�/�TDc@��5�K��q4�G<9ǡ|0�|cɧb<����Р���F�#|<X!s���S�u�>�{��t�S��_Q�
Я����k_�JBST$)KM�L��)�J0
���"t�KB"�du��'BթI�E���[o����cP�۱���n��c
-
���+�D�E