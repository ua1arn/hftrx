��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^�u��]]��c���Nd�e�@Ѱ��iw6���=uC�Q�׾���VL�����EQ<gS�Jdq���<��;^�<[0HFI�W�W05��p*x��$���[��l]/�a�a�U���k�bS���c���;d�#�{7H�2ŋ��J�3��Gqn(Q�¡l��uw��:GV|����J�'[MU��0qZ!��*T�P6٫g"���(�4s�4�f���_���3���=�3|�7�(�n¶Ē��P��ٺRd�Pa��vH�r];4�\w����F�XX��Q�AF%\�#�eM�5�K�5˧־}�G�s���P����a�[�gƉ��銴6	I���&|*�g�(���`|�G�d�q�jz��2��I1 ����׼ܲ�5FZc��V��\�ee�!�"�ĉ."�,�� 5�ݕ�?C�P��{З�wPt*��@ܯ����g�/����u��N��1P!�F��R��U��\|z���;5���d���Ȓ�w�}B��5�z�M�����+S�!�
��$�36%�f��Q�\�b�Jr;�Gn��Ng��6,י�����>9�x.r��u�3vڠ��M���/�f�s`�g����J�9$��6UGV!�ʟ�7�3L긚	*�����i�5T�rY�I���G�ϐ\�[���ᄯ81��vN�	�I�\	��W吟C�!�OQǳ��Ҹ�?��_���蚡�違h��v�|�v�E��n��=�������ڏ��ma.��<݂_�����y\b�V��p�f���E���>8� �t+�x"�ݷ/�]��6?�>"I�R���u�0�����%kĵ���`¤	������e���M�aXy�z����HbG�	������,B��M�G��]�d�X}��H�l��n sPt>����^t�����'^&�.�`XQ�)]�qX8O����O;��EN�����O�"�GCu�XLQ+`Bow�;f5�m �?#n��.EV^���#�>?�C�����̼�}���j~�����KC��W��S��8m��m��V��_�L�o��@Q�wq4ٛ5A4�Y[��YWm���#��������~��4%�v�6ܵ�}!>��(:�F>��ډ[��jLVN������$��n?m���A79���~�@���4s�HD�@߯�����`b�UU˭dj��l5��yECY��G��S�Ѫ_I�8�����Tn��}b��r+��#��E�S�G�s�Nt�1�p7�v%b��ݾ�;A�rŻ@��Yj�-%B���P�Þ\m�������9�wdTHo�)�	� ������&_3�oN��9j��Q|����#1� < _yc�U�x9ZFB>��\���}�q�`y�69iC*Pܩ�(X>q�s��O����Ln���9|��z9��:�u A�+� ~ȅ1��uy^4YHۋ�����4廥�J�?����x������j0x��]@�$��"������:g��t��:9\/���Pn�^$ aQ=xZrj;׼�1pi�Ǝ=Zb� ��JKq�̦�D��^Z�x��V��)��{<�H�Qa��L@���v�浽��o��Mf9U�||�9h
�?D���P����-S��)j*�v'iiP���ej��8�GX�y��ig%I횑�1�m�&��Jfue�a{ڞ-.f��ɇ��OY�WP�g�	�5Ёo��YM�e�Y�����%A 1d��c�#{�g:*} ��7�I\*�����P2R�e��7��*p��أ~�'��w���9��j�^X����Y�#CϿ<z�m�s�ǿ�����'��v��#r1��~�����e�o8����-<�~Z��Аj<F͠%F��]���n��*��;�ByC���9Ȋ��j�c`@
�OR͟�������J��љ]��[�+3�֚cϬ�ǜ?[�+%�rd�ԡ��N��zf�� �ܮ��
i���r���Z�=��w�?="I���tdQ�E�p�\�.�FB�%P>M�����#;�	E g�x�M�p�����;�܊��i�E��I�Iǆ�ɥǫ��8V�����$6�Y�5�������]@{s���Yu"}�2�d�_�}9�pf�?g�&G�Dں\EW�p�B
>�o��CU������Π{Ĉ�M����ĬE�{�q�I��"܂]5������>���̡gZ��J��Zna'�Ћ�p�vʨ��꫎�k��ŋ�5�,��q�oP�� aWQ�Ev�jz^B�kk�KN<�K�W�ީY�	qb�Ǯ:�}��� \G�z�{� c����ƥc�N�� � H�)�<F�sK����Yo�sUn}�E�'���4T�`1B+��<��^���۠��>D��b��#��*�h�5�T�s=�B����R��	N" 'p6M��̰�wGq�����\3�	��SYf������
�;Z�%��\0yB<1ߊ���H���;G�^ƎE��������㞰����[Q�^e���/����Na�o[�&X� ��e��W��M�,��E�x�BWA�#�����2)m*\9~�5��"���sH��Rv���^��k�ˤz��1w�63e׈�8��sU��^NңZ�-�<��u���'�y��2�Cx�`�0J��#gZ�w��@o��@.��`^.�WzZj��$��0mP�:��#e�:����ٚU�d�G�����Io(˫(���s��x՟t�[L���d��*b��.h_?�4;�y	#����>���b#�v��[�I~�?��ꐧ�*'	�H��,��)@��U�]Y��:t��4ȬX@��T;Q�Y����_�IrC{sVmrv�����;�Yi7Fb�nx(sÌv�C�U����C�h��y�Nl�������ۋF� H���gU�%Q>�d��Qݱ����w�a�h�\�|�=�ZΊ���Մ�w�6�lI,�"�j6��n{�V�uvQ]�Y���gɨ�6Í��-�x)�nf�c���}|���.L�$�	�I�톐6�%��� U_�qf�����2 GjR~�!��3��ҩ�Ԓt��u	�O��,Ɯ�?i�%��
�T]�����~��t�a^2̖|��ESL�>�����ѬL��BQ�-�':3�b �x�wG_��:j-+eYk�@�6��9�D1p;�,��8�[�\�K_�N�a7TЦz��S��iEu�Ğ3���Ҥ(�~�^�C|�]��?��2v�j��Y6̦({6�Gӂ5[7B�.;FsG��*B���;z�8�9���s�*)�xŽ͹��4��T<�
�-q�T
��[�4��t���*�c�lG�@���q.��$t-7��p�WOf��w$�v%vO�~�����pyu���Y@��W]px��s����-�[](���^�T7
�7�y%����Le*"�Cl���6d!NB�>�ߑ������D�*�f����b�:Lz?����I��ڱ$����t�ϧ����|��߈z��nF��:J�>o\ ꇃ�n�i����[ޑ��:(x��n��KmH�N2f�������lIw���(��Zn���V!k&.'�Ѻ�+��)h��0�H[��7�VU�����]�&�W���t���@N�}��q���<?��#P�y:�fSb8���:t/l���U	�אѤ���!jđ=��������־�A]�C~q�b�OR|����㛅���j�/�M��K{]�o�I,'g��t%�uA��Ҏ(./��L� �u~�"_��7j�yp�>�ϥ�'����ڸt=�D�M'R�+��<�O�8�M�����e璿���_�1�ˉy>Gh��σ����o�ܞLZ���;���ye�0B�8�`J��	v�������jO?+���$?�����Bqs0��	��Am	���^�t	j�W�� �Nj��V�P{,-rӤ|��)��*r�Q�2��ͤT���O��y�V�E�o���(h}I���vЬ�6��o�F�S��e��Ǥ����<:�_��_�c���-<�C�r��F����3A�v�A�UT��tp_��l�n�=p6��BT�$�Raa���!th�g�+mB�O1�7���Z�|�2���	K�!r�z�b�̰[^i*�y��̻�%�D�s�+�iy�/e�+�8gJ�7�2t,�f0͸~��Ĉ��0��vt�X?йjd,���[G�����O� `�T��PO�tV��,L�6��jg�|���E�XE�|:4a؇WݹvV�Qw��U�����
N��_p^c*�n���f�{qC�a�O���n��!���[�k�T�1�0�_+�η�'-3�R�c�i�{�R	�����E���_F!}ǎ��^�'Đ6,��z@r@����|'�x�;��'�D ��Q��y�_b�����vX�H�]��`쫹��e�~��O��9b��Z�W=�@8?�Zj��yc��Sh�}h���B�S.�{5)z;�1��'	��(T�y\�J��ډ����d�z�&Q�Z���"oX@�����C���F�LА�^%;E}�Rf����Yk
D�6U�R`�|YKw�����u�_W�f�TZI�N8q�J�U�Im-^�͜j��Z�~U�
�����ۘ�*��U��u�4�ˌ��(�m��?A.�����+�ݕ⌈p[gX�HeDR/R����h�R(,���N�m'{�e���q ��K������L�/[�Jk��,UM�DKo���>Np���r���+YĖ��߇t�n�8,�Ɯr�7��d�k̑s�_������Yc,��+���{H��^����->\�Ә����S�4���XH�5V����ģjX�	.�Ҟo�Dr菉�B.ïv�U�V�Q?�7���AL�w���m���� ���E��}af�_��tj"��{�Ӑ���B�ѫ���.;pLu�7�B�CΞ�^o��3�$ ���se��.����qY� �p���Z�fl�U�#�����N�>A�%�\��ȹ��i�#�����˄}�1~�$����6?� p��Р�
l��g;s�h�`�m�	�rQJ"^���TK�����㨻q�/*"�$�-²>a�g���<?2���*ْ��I�����(w9� �"�he����fBƺ�J���̿_�VJ`/��Ƥ�	rN�}8#��&o��٣}��@,gu]�A�S�J��s���{����K.�������6���.�?j"/�~(2����W+J��::�	���W�	E����װT	�p=B��r�����O��� ��e'�5GfZ�����x8O��nSdG��1�'p� MYo��?�@4���W�Kޤ?{[g1̝�Э%z��p!���_�r�1C���:�D�J�^��.j6���[by)���;�u;��[�Y�ڰ���$9��ī8ρ�B`�{�ӛ���
S�����Nf�N�[�i�������d���^?�J��Z\d<�@=��n�����h(���Ɣ�jN��	��+����9J�8	����!x#��Z�I�W7�ey��T�����ׅޢ������"�*�@>��O%��Go��=oꗱ�ŗi~O��}�<s�_��2>�^>�<��߆�Z9��"��HKKK���ɒxU@H�6����GXv5�w�z��*��Yz�.�0���43��y��8�j_�e�����d?e����:ޏta��� �u���T�Zy�Œ:v�X�N���r8���~*�dfdXY2���N#���Cb0gi\���j�������k��C�L��U�\�: F�8e*WҦ�n�q��.��F��Y�Pբ�J���u�>�B8Jao��8g���P��Z;�.���?������h����U����I�{b�P�k|��6�.5���F�|�jw�˅��gyv�SGQ���(��u�}~����!�';w+���	&K9���j3��'�#?3��
b����\G�"��r���.��� �[è'�/�?��?���O��'~���yd����T�FM��N)�%	w�ڏ�T�o����X���Vs��xY�rt�>�\$����S���Q�EV�ig��-��������|��5��ף��<"@�\ 'M�A�Nb��¶�Z��8��N�%����=}ߊ��y<����K�J�̐$��?s<�7���t�ȃ8{{XK�+W+]cD?0YE��E�)������շ�BJ �U:M�LB����q�GXg8�|U`\%K�/��J=
��;�k�a�I��N����qK5�w�NsE.N3�)��'�����߫P�;�O^���8�Qʆ�l%�ð��������T����кn�+��T|��*�) J�R�=�G�w$���2��3d-#x�eW�{�5r�c�e���>f����;�9�el�[�X������R���e�%n](���{t����5Aai�]d`�%��Jy]e�VViM��˒)�@f�#�e�ױ��K8�Ehg�-���
�x0�۝D�13�������[�p��dn��&��d�<�6����n�� ���uJ@(�&T|ې�}�O���j5*�昽}�&b�G<�K��g���_F1�Vp�2�h\��U���5�Z,_Y����n�+y��d~K�+}</�S�L�b�
�}��=�����տV�M�A��<�\oJ�f�׌=�oC-��
��&�Ɓ�Y}�*��y}o�0v���98sV��N25���@�7y�9[K��XH����c������~�*���@�8FV^`����`u�������śr��;lĦ�_�!��n$�9��
_SN��"�^�� qR�����R�<N
�KZw�K���(>������ͼ;��绐Z��>�N�"H3f��.R���߰���Ē�'����e;;��% S�^��x�b����U\v#��x�QS;��U�����t�$h�3p_"�RH0���c��z��ܰ�e�O�Vϑg
 �cR� 4z��Iꛫ�,����ir$ܔᎉ�E��q�݀p��������U�ʇ��%/��az}��b� -�h�����OwV��=�	��dU+��@ "��&��>�<��j�yN���1��1EzFeu7�bI=��ڢ��ւs�X/��`{c�pjx}hߊ��A�L�k�i���1�N�D�rt�X��Y�fRG�U��d�A���K�}�[F5:���V�(:	ZXҌi�a�O�M�I��I�Uρ�[�0[���W;W�cu�AR�벰p��̻�����+���Q68sM���2���j���9r�w��Z�v
uIR|OjA��+���Gq442x/QAm��>�D\�$�3[7̋�KR���g��2�_5�w�«�j�=2*`9���g�����z�M�����9Dt���/z���������}
8"���
��	�Z���%��<d�E��5Oʐ�@��� �`b������_��v��C.��<��b�M�M��Iq�����պ�R�����k�>�]���B�+��`������4=�5Y�#.k��K��+K�fT����&�ޞ�Y�H]�����s�8��"{a��_�v�L�������57��ED?�F�K�V�O�^�M"F�ki��i�s���=`9��oU�L�r$f�>�E�����]��?mm����cO`��	:�{�bF��0����ъc@j�]��.�u��F�<(����#j�xL�Y&o5(��O-;[F�Їp��pDPޒ8ӿ�Q2�Q����c;�D�GV��X���%�-`�����MҾvX�eM_�!1�H2�3�b�ލĠZ�Cٵ�Y��N[���2 �`��lTmh5?[��n��M� g&���7�cS���~I +�vX(q�o�_M-'�k���a�6�ĳ�+ÃϾ9$q�����RB��@��A�Q�q�Jb���.<92Fd�Z�d_Eu��`B&t���7�LS�� >�[G �9�\x�G���h�Ȅ�b���dh���N�)�Rn}o&�e���L�C�0H�����q��~�n�skG���'\{�l<�T�.D�)I���r�@/�K奊��n�:/�_9�0*��L���A]�Gz57���С�m@LJ
�v^�����>D<��b���Ӄ͠>T��aϗu_�O�B��2�FH�y	�#�k0]�S`�i��݈]v������}S��bɞ,�8R��}�K<�e:�'�)�5�>F�^xX������#��I'�"��y#\ �2,L����V��Z8�CMU��3�\W�gS>K��ХRG�q�G�?�7[��b���m��~�ȰXW#��q��P�1up����:�i�OFr�2n����HU�KUy5Ԡ�% X"����N�C\��]���d�-|W�:&8�Y��N� �T>ˮ��4�Z����=
	�p��{�=�7�v��C����y-�(]<S��	��NT4�|b�F�Ůc�b�H,?�|C�ɀ�ř̆���ݥ�S��;�=�r�Ǜ��l�?�����]Qb����} k����5#"�u��z����u͉�*�w�id��H�a�ZGƅ����2��i��R8cy�Y��S�zb)4�CJ�B'KM�X�����F�)Д�p�Ԥ�+��)綦��f��ׂC��1��<�a\3�&M�(��!���`k����gж�v�!� �� �]b���V�h�*	{����s�³�|�J%�h�br�Iz�U.�h���=o(h���}ݤ3��t�*R\^�.��1������\���oү�xdƷ�cٱ��Jr�Z���:߇��_���kEN\��~cՂ� e�go`�'���v�S�ߚ{��|�g�*�k^|��^ߑ��VM{:T,:�j��;���S�+]�
)ϡ7S�*��d��.����w�m���;�k�H� P�a���iލTK����03:�G�r��V���\�����k��PJf�6``�D6}��A�FK�M��ݻr��*�.u�'�I��Z,��Y��e��Ȭ)���U��N�c;��M2^�Fq��~���$.��θW�I��y�׻�4f���Cb�"��r[j�$Y��f�,��� �W���mC��G]t���X8[�����`�ʼ����EH2��4���h�m����������YT��l��O6�lڟ�+�M������UcTDE��/�B�e��<<��`8q��t�����kHc�82P:���x�!��t����Jw,%*B�̬ �V����n��h^:hH �+^�vk�� ��t���j@�L/�6����T�A5�L)��e�xoI�����f�D�B���}��"GhUeQ��t�	�'��;�##5�X�dzX䫕(�U��J���.8".bi�l������m���jOn��Ҧ�#g���M���yK�ès��.+�wNXh5'J[��`čXk�;��u2u�E�F�q���Uh���Փ��E�dD?�C��* C��c��N,~\w}N"B6��Vel� �� <e���S^1��I����צˠ~@eK��矇��u�uW\!��*��C&&�L=?s���*P3�"����-뀠�ˀ�p]~zk���R�� ���[�O K���4�LgW=D��{J��p�88]��	(�-�<���u�W���kJ�� �0:���'���Lp�	��Y��T$��e>��bE�P��������$Sa%B�ՍrB��ڃ�o׷yD#�G�Z����U�^=^꿴5gO�ۉhQ���wzJQV�𦇃��������!c��qP9\J��	f�a��ց�����z�
�%��30��߻@�)B(SR�o������0�L]7Ɋ���a�j�zdb��a��-�����&�ѧ�������V��ꢕ=�{QB�p<Ifgѫ�yn�	]�E��	� Ȃ
�d�j������-�3P�2�X�r'͓<rsBS`TJa�2�Iy(��,����P�o�S�ux
ӫ����u�"�����O�(=M]�zc�<��%X�=��ئ�U�U�O�t���q��8*��"�y��%�D,��>b����8w����� �0`K���[@j���Z�1�����q_QpJ�O�a��oݢs�
�ٚ�������c��(AiӜmWB��q`��)���ݍB�7M|��7]������?6u�m��^��vL��/@kL5zv��w��b��52`�%����S"���px�œ�O�J6��h�W�;+�\�2�����ZQ.�tig�˼��y ��1g�S 溼@°u���п�O�W�����dZ�U��u�� �Bߊ��L�q��dj��A�ĺN����e�a%��}t��^#�0K9�"����3���"s֎�ƃM���A���-�����U905{���k|?��ޭ�@~�=w^1o3����'ɣBk�F��/�>�c���
�4��Bu�=8-m�܋��̎S�lEWW�>M�1&���;Y��\x��pH9N�4ڰn���,Ш݆��E-H,؂ಃ�(�D�ȸ��E��O^~�#�3D�VH+	ak��l��N�yQ���׎;^5g��f{e#j��Bz���|-B����mA���#���+�_�GK(�1H�����Jd���S��6��s6;i�l��&����Yp��R9���kX!�V#A�%q?�i����+��om��_��Y�Fy�cFaQ�l!�$�ⴛ�LzsL�{�^Z�T9!�b
).���c�?*v&���8�]P���l9�������oq��.t�k`d��Co��q ��%�E�8�+�`��aid�С��v�g/}�4E~�GTI��]h/8r�U꿦� ��)���￥�\�	}�r��,`�PQC�YQ`)��%�����w%=�D�uy�y��Iu�ݹK"�×�����g4SD����cE�J��Z���цB̲z ȅ�ǅx���ҋ _�+�{� �;�͞άmhi�=�a�3�1lIy����1�I�^���3�D�Vw�0�������b�0�#&��x����h�֖>O�ⷅH$�կ(�Hcd��mw-������`���퉘��Xqy$2���*��U����&�3Α��W_M�pf �Ő ��H��1�}�7���W�1����|��Z�6QT�\G�Dr�	p���
J�@W����H׏g��a��H��xxs�?�����s�7Ń�w�
f�'ԝ@.b��h�<s_�V��CK����5���z�� �?���x_��Ր�`���qG����'>�:���`���B��h-&��?E�m.��uf��Vr��N|v�������tY7s�����#��A�?#7�i#�a�m���,����DU���������֯�\R�\��[��΍"�>5���0in�p�5�;5�V{kŚ���VS�5����(��-4\�䊜���9���畃�"/Cj	*g4���0p�'i�����e�M9[��@s��ؤ:�4��iZ�I�>S�C4�z�p3k��;�?(,;����deХ�zfD��!�g����W�㔵�(*�~�Mfuc�+v�p�)'6�+��w��O��a��������.�K{��п��|��~R7������;/*��%�>R	S����|Cײ�t �B��M�����ƕ�_�`���*
P� #�vb�I�#�\#�I�0���q�����qp��������`� t�7
��$��#x�جL>KS���u�w������a#N8��]���'r$e��劉��/�����-7�f���*�A��ZB߫�J�S���-g'���)�N�
"m(ގ�|M]��č��y;i�Ӕc�/�� _^q�"��0i����@׫ٗi��u�
�jA5�7���0��d�l���귮�7��V�h��,Sb>���i��f��k�x�3��N?���r n2��S�l�]2���M��x2�	+�hi�x���8+sBy�x�O�{�~�_�:R��\C��;7А�����Շ�3�y��d��.4W/��{�]��uR�2�7~�w�h�� ���e��9Cݞ-G��2�d	@�jǤ�.�p�eK�q���ُ�Ȱ���:�>�e�HƐ_bmza8 Qty��RH�)1,<(e0����I)�|��y�i�EMwP������/�#`�τ�L$�bIS�_�P6�R�x��*o��zǴ�1�db�-:<V$#-��L�J�o�ͮ|�/���۟7�F>�	��͛_�~�o��u��l`9�O#0��Ν������b��y�Y����G�Q��qFF����ʋt2䯫J?П���a�	|g*�#O���/�� �v�	�0mRq���!�gQ�Y���o�|����,�9OT���Ȣh�Z����J:�zh(�a�5t{���(��,��B{ 
��C3=@*%�[R��
Y|��0
�����U�v�0�T�p�Y�݆��r����Ǉ@
ϗ��暿k��{�fؘB�`wn佁�`�!,��w�7jXa�@$�|q<��8��Wܬ �Yŕ��7g��uq������]�u
��Υњ�0���
$�_<U���ժ9��r����:F�/����|�i�3<wy�}�6�o�M�0�Fk���f:�Q��)`�~�d�;>pu�/)K9��r��y��Y��F�4.�`�?	 ���#�ҿv ���O�-��;K�`z�q��0�n�%L�^�?&mDeR|%ŗt����_�yU`c-��ړ�[��X�s,��œv�����`w�H�4����Y�}Z?�e���j�|�H���&quJ�Я���U���(��0���$]�rĿI2��4FuG߈Y�mh��ؑ�'@+$�сJ�z��`ż06!4�������(;k[D�:�Y�y�-��V���;�8%A����So����Ia���\���[+kԧ�j]A���=ˍ�̱�e��ބ��Π�2d�H�q��IPS
}�X��ݮċ��M*�|��@&��T����r
�G9�VȚu���!�P�Os(�E��64�F��P:��K��C8��٫ %����l���Q��3�"�`4F�g3$�=���v@]�A|2R{s������tzt6���+=W��y�C�#2�����Q^�Ə4����5����%���tv�i�����J3�$��E}��6bIt���i��A�E��UJu�n����#��b�Z�.�hH>}�Ϩ���L���L��=���`B�.�Wj\}�:�U6��L#�����`� �O���~v�e���|oH�(����º�߸Q�}cB����!@���n��9BO���/Ka���ʹ�l�:e�eT���w��[ [�v�07�KۤI!�Ɯw�L�)����ow�V���g3Aճh4^e���g����m��˒��WO��?�8�;����R��}�8�.�~Oz%`?J����QG). ��0�is��$�lu۸����(y�a��HHƺ�%�>�a��o�!�,��9{"_0��jyK�8;��^#���0/�]?2EB3���n�4/'�°��li�F<��E�ϭ�"Oŋ?�[��/���A���d�;�����'����T�!��{A{ �'�n}O:�Dm/�p+$Dp�t/�q�B��F��X��&�v��ABs)�ې�t���U�I{Aգ���u9*�U����~���q��Qr����|�5�y�"�-����H�u
[z�\�D��i}�m�����8��HU~�xm<���U|c܎ܴ���'j:���ˍ�
�)�Մt��7,.���?�����0�H�DSuk�{<���,���7#[�U�W����ģpp\��?�\�oi�3e���5*����v%4�EK���p��� �M<�}���j7�bN��'�g�r}BH�]#�7�fr�E��ߓ�w#Q#�)�ר���a��u��F'6#�&�Q�ƶ)t�_�R���"��d�GfižH�h!����;�e�Ǻv�,L��f�;=̱�U����;p{i���9�[��-N�q� V�U�"!q�t!CX���2]�$)Qޤp�Z#�q+�bܩ�:�)aR`vձ"�^�h��@����	�3���O��c�1*��*�=1�\TI3�V4~��^��=�4�j�;e^2�YyS��n-�'����T"?.�YT�3�eGszf��&ˡ�WH�ytzx�����-�%��iR|���S��C�3��ږ�~��ԃ�ngb.���E�u=���/c���/��q!�R��d��}��l��8�R2Gߨo�Ǒ�T�N�B��!˰�Me�K�H���iX�v�rÊpУ�.,���!�2���'týY+2����T�F���I4��Pe�Y��Vj�����n���
L�I��O�傎3fG�^|��փ����c{H�<u�$Y����.�?{��>�ԇ���㦀W���}O�$j�B0p�j���axg��/�U^߇�M`(43/��\�#�z^�R�<o �<L��	��L!�A'w��ŵ��*��[W��7�����VY*�AsW#��ӗ��c�5��LFh!L+?�c���QcUΡ*dr0\R���.�E�����{΃Pi͛�Lڷ�F�B���{��K��Gtd�_�؞�!�-X@�/J[��ew��E�XCXv`cJ�X�l�TK�W�h���߽��cC,�@�ۑ�&<2�����'�s�*J����.�O��j)��]�+�ZE-Odh���H�ި���w�T]Cw�P1�����#!��/��+��;B�}�؅'�����~�ir�lYD�(�,��8��p�����;S-h��ʃ�[��K+�CUkx�3֔3�z����>2�mSj��H�#��h��6U݇H>'�A�`��Y�}>%�Y�$�U�%f	~�}��}�Gz1��6Vц�E̠�C��O�iL�݁v�d���(I�Ni��wy��|�g����\ChE���.)Rfx����lŒ{dls�v�tź�|Vexx��,e�U��)�q� �l��sl�D�K����j#_��_]"�����e}�HP�L�E,�ӿ�š��k��O���VEgR�}���\��֯oZ���S!��I�E;�@�a���-�r��/(R��f��$©n�t�JQ�T7f����msO�2��1�%4n�]�+n�h���ΪR�l�o�,{>sdaD��G�WĊ+[�C=y��1�jл=�J�[0O�:-k�����Z:�L<`qbqk�H�d�ɓ6�P�k0|k�"��A�<���k<���-DF#SAJ�������FS*�Ն�|A�����%)r�o1��*ɡ�{�����Q��Ӓ�o�F����aM�e���
ՒkϞ"A�w��>��Jk+��m
1��;yw�J�B����&%��A �Z�|�l�jb�?�Q�$��~=c�|�/J���W~��"4��k0�� j$8�~K̪��s���H�Z6ZmH6��mG��e%��f�
�����\�G��{��;q�k^z��a/Q��x��o�(~e��@n��~Iʌt�6�����@&���%p��槖BCn����F�T��,P��5T��9�";F�^Jɩ�4B��H���s�E�����Lk�+
��Z6��/���Ej����4iy�A����N��ox�b���`,����Α���'��Y�p�W-P� zbu�[�V���,�����y��^8Mď�ybh�Cg�E\��oF|�2��屨�kIi�����$0�J�ul�c�Qd��ܭ-�!ϒ�P-��f��;�PT ��X��6���_�CE�s%���88��f%GB[��~��_f�&'Ӳv��+� ��<��n�%�����n��"�����Q���kV�[ rDth����(2�
gKbܛ	ٻBΩ� =x6�̴s�,�j��2��][�k)>%sP,�[.>B��.;N�D��b����Vs9,�*�?������M�R���L��@��Ot��2�\濫��q�	��V��0��\oH�0Ey�ڻ��WVHO�� ��˛�dA~���sE��i2��t&���Cxr�YfqC���F�r��L"a^�,�|�����h�a�z�f�8����1��(3M���o| oJ��������'���3�
�X-�6w	`Լ|�~�*�;)fn:HgM�5L�6r,��?��!������ξ��?�u�i��ȕ��neݹ�:pqz
��N�9bs�G}�b������L�y��qR�7*�nO�D��Tp��T��Fz�l���I�}>l���]�C61��Ozc, E����r(C�Ӻr��u5�e����_Tc4n�-��B.���gC�k����`'�q�ɪ3:u��X�U�hݥ� ��֏�Og�k#댩�$��@^��CVh��)�Qhf=)	?ρ�,^Ú���T�R��1ff������ٞ��z[�˗9��}�2?��I�D}��x�Ԁ�H셤8e� ��Ω�΋����e���s��c��nA�ѫ��k)w�d/�	m�Y�� Ce�pE���q;g��1�l��9L7T)�]�d"d$�0%��n�U(��p4c`��=��p���#�l�T��&O�*g�d�"��8��
I590���itH!NK���ZS�~-;�T`q���ۄs��^�s�CA�`���B��|�����(Y��"����s���lvjiR {Æ����V�}{���%�^C�jyC+-���܀D����Ze�:�D@B�����A�"��<�Lk횫yez�SJ�oC�+��M�y�F4�I�����G\C��h��T� i��$�:c@�EYkȈo�˞m<u�|�*ދv�s�A��0�I�zy����sc�pX�>�!�GbQ������@HX}o���m���w!