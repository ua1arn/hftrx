��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga���<�\��J�ιϛ�������tFpF�)���u-�6k
���AY�vݥ�WpD��G5��������cF$`�� ˄�.�蒡�q83de��+'d����ĳ.�L�8& �q��V[��p9KY����!�ۊńR���w�q�����k�M���`���
bċ�T�y���$�Y�H<�(�u`�>��˼����̆�i�]�/�<�a-�^)qYOA�èMX?��_��d�akN����NT�(�&k����׈F�ĠG�JA��)Oo���6n�ne�ƾ�D@��>��l]����]ś/���䁌��� n]�"�6��N3)h�@�b�U*L��r[��eK���`x�)�$c5z�o���2շp�hO-Do����e%��������!OoK���)�4��[w�(6V���Fd�:w� 33���y��/Ng�rHW<�Щ�~Yx3>t������c��A��xK�J�c�'�Xi�G�6J�:'c"q��-�]%�T�4�Hr�Ge�gejm��y���V����U�<5OT30����Y@�S�X�qcxj�J�#~����� c�-�x�z����>�|!��dm��!���|J��͛Nݸ9�R����j��v�٫��0]}
o��x;
PN�Z�p]�]#˧ͪ��mes�S���}��Q0fW�K�s�	Uto�I�sj�C�u����2�sx��=�����T�[���u��3;m�"��T>�s���d0Z��"ԍ���I�o�y����"-ǝ�MT�N���v��q��'����z��A"�Q��3�n'*�{��K�F�/���1H4�$i��b��������B��O|WQ�	�����vA8���L��?k���3�� %�H.Z輄��HG���6�܋�ꚉ^p'��e2�7H��7�d�VG����L��iA���cz��á�Y�tf�oo٦�2hB�M���keɕ�9��K��L$]	eD��PZ�yhhplD^��W��6ѱ������| /�7M��vݵ�e�e�C'p�k���J�;a������Z|�40w^�o�<:u0߽H�؎�`��� �i�bqnƭ��=<m��{��דIߖ�..Ml�>�W�g��092�G�^���H 1X:$2�a�]�v�
j
�x�����k�L�
*�P4:�!�m+Yv�A1?��5r�@f�~�B/$,]S�)t�����_��[f�	�55F�J��Y���1�lWB4���T�r�bHs��h�؂́�h�rO<��������v��	j͸>�J�=�pH��@5�\�KM��'B��0&}6ߪ���ZƼ&��̴��
��E�7斦.�̏�� 7���~`fa�*��S��=�
goCN����f9j�{�M�74��!�B�~b�
ȸ;���ʣ$� �hx9'L�݆��g�ۚ�e��߈����l��Rn�J󂄭���{4��gA2� �q��p/	�ϱ2?
�D@��E�(8��n��:v�v� ��v��<���)vѧ���"��{FM�bR�53����2�8m`v�"�P��c��5]���F$�Qz�{�ۀ��`KWD�w�2�1yXE�S��P�&�����!���v��W�t&�\C��1�d����-M]ę ~G�p��-UP7��B��ͯss"GL+F|�R� ��VA��ط�M�Z�/��EВ�o��(A|L��E,�����N��F��/ݽi��"�B�L3�(6D[�}��)����`nGĹ�5�"�
��e�C�%��2�k`v� :7:�?T�l{���!���Cޞ�s�|9�]��n��QA��s7�V�y(���`%�>��l�A95��Ԃ&K��6N�	.��:_`�Ɨ��F��k!���B�pȧ
�߃�xr|����CR�Ȇ8�z�̖��H�vJ�
���u�B&��1�g�L���������9�Vp�,�~��y�H�ʲ�%�v%�V��L,��`�y���q�_�˰����Mf�:S�%Vxg�֋��?�v����󄣟n��K/BH���" �rg�>KXد7�b�8�!w�E��_!����\F ~x�:���А06�[�u1�j¨6v��,���B=f�ə���o>Y�n��nDM& LI�R6U�mۛ�I4�,�Y�hs	�u@$�Ll��M�B-E$��M��9�^��N4k���c�����X������n�X�Y���(�;#,+�K�~5�JЗ�y8^���x�dB�8�^O_��? q�K(�ӧnZ�򳳢c5��`'����Oّ�+3ii�P.4�R�Hp�@[�
�hz��Þy:��ʓ}%LNO�tID�����q��hF�=B!I�=	?#�4oH���X�45�\l��h��eAQ	fv�[�U���΃��ܪ�E��d.�첈��\]Z:��X�M�c=frs������]m���g`aյj�zH��(@U	�$
�Y���o�W�J�Y�X���Y� �J4�1mu��(��v�KϢ��M9d��hvH�3�U	��� %�\q7��o��%	=	psL��ɺ��j�	OV�{�8�=�,j���oVk�Θ�iW1��lch��(�2%|�5N~��l�U�M����{V��[�F��3f� �
�T�	|��"8���f��'���z<	g�rL����G����"��U�\��E��*�I$���D�bފ��p��%,ݝ$_+�/��S����J�9��	kp��ί}�,.���xU�F���:�Q(��e��X�5FfyUM�v��N���!!*k� g��>X��t�a��FaS�Ἂ<�,��l��(z�X[f%N�|��Y���� ��Z�:D��S� :�fK���v-dy���ܟ���EAa�ՔDr��Թf^��8��Lz��"�"��:>#u����O@ �g�[Y�P�X���+��qO�*Ww�Nl«�)7ð����aw~���V�Ε����-�k��"�L���K.��*m���0lo~�Co���߫�Y� ;]��3�F�y�	��}�>�L��!�,Q���~�d�`�?A����L���D��t|�ޥz�����J�O��W�� ����[��v5�j��7o�z�:g��z�[U;����/���=����j1@
mb�b�_+�W��%S��܇��3�;�9�����[ղf�0 �1�y��0�GD~�r��aSz�8M��*�:�z �C�w���>�$��Ta|����]�[��D�'��J�$��:�,��vٜ��C7P2Ar��Gw��D���Ic4���EG�~�tT���\�y$"�WY��?C�D r�ƭ*��M��Ȕ'a�/���=6��C��Cˬ{O��h*����}�����۞���,�߆�~!'�O�~�����������%��I���։����/b	�n�!uk	��;}5������:����ڙ䏎:�����ۀpi[�'�鑁�,��P�ɵU�s`�%0�a����U]D�����b���������,�*O�,�U�L����?M��� Kr勚A���i�M�n�(�!�N�{vEC��a<�:�l�ӏ��.� :1��Ip	�󠳚��H�:Y���s���AF�V`[�A7zׂ�IBV'�G�uh�A�nH�Dʗ�����'�\՗W���;��oIV���k���Rz�m	�j˕n����xр�w�bƏ9���e-"_dpl���=%��5�2&���{xL]��L�ڂAq�:�$��b�����Kp'gv�B�ua�yf��F����|\O}w`s~z�x)L�eo��f(�_$~ϴ�����z�1��g��R���oxN����o��2��\ ���]ŕ%���.�/Fv���	8�����to�/��S��J�������w���a��T�wZ��L�}����P�v�z*�o����K�����FsW듟퀯�$@�0,1U�M��wE4�#�48U�֪�ȖX�}�m?r�Yߖ���Fi���7Ⱑ�-|6boX	�)�L��Ir9jm�ø��)���3�Ɣ�^�����3�����U	�%�9���|�諏�[53��)���{Tk,/m�%D�y��4�}AQ�8�gT/(W�X1{%�dD��_ys X~P�ĺ�2@��t��}{�+���R��u:���ݶvPP��� +p�P�x�PL{��m��D	�!�J����"#5�5����ZӥU���o]�74�F�Or!lt}3=�l��A`��q�����ڐ�*7w�`��h�J�z��i�@��᰾@	q���5��f4Q�y9������,*"�Ml�|�Ұ���r�@p`��P�gp){x;հ `�.}��E9�S:��蚤Tn��L�s oā��(8H�:8�k��撉���%U�{���2��JvJ[q�U�ba��Gh��h��o!�%��"��$9$�o�|�&�|�<�����/�ۮ�©/{�j�@-��A[� �b,_�4p���~�b�H9�4�9L�P./T�G�+/B�� 0�9�����\�/�LB���K%������h� XE�7�9(v/����G
��F��M�b%�V5dK^�栃�bΈ�6�2���q/�� �<� :���-�ɋL�D��6��P�13-4����6`��M�'�O�����7�<�'�A)6Q��@��A�Y�G��jt8p���Sg%	���x���!m���9vREH�����n�Xb�B ѽ�^���تx���Cp<�$�ʋ�l�7;9�m��z��w�(
ݱ����7q^�|��CƪH�°�3�yȓ��y8� *�/=� ��!I[��Ӛ����ˋCg�������ݡuW�G��K��4t��C-��']����w���Jh�����7���|숐��@!�k���A�?����J�nX7��������4$쑌��zV#=����G�w�t@[�m7�t18\�����<�%��\�eR���g���g�?�V���\uP���A^U����*���Z;��?��K柵3�����)�/2�&�@��4��֓U�=*x�6"�	�U�0��Et��] �Av���pQt0��ht#8�ze�'���j�%���E�t�P��#�w��Ci6����^��
��x00�D����.2C��}�u��F礆KY�rߓqn���)�:��&�'�i��f��\*_�c�i�����S/�&Ѓ���`�:�(\'^T���,G>w�{k�}���n���ZZ2Q����Dd�P�Ƚ�	��Ϣ�EJ��柯��͊P��3D'�k9�b���SN����YvArZ��1<͇���;ޯ�0�l���y��U��Af*ğQ�q��+R���>L�d�{+�h1s�0�a��Q�A�}if��X~�|*�Ѹ'�o�aoͪ��qwa��f� �͗y�i=���}���[�ױ('b�d�d�1�Qa��h=�Y��=)�e��ϙ��Z�6J	x6��J��&7
5�#
���9�l<"�hy�7�o�ۜ�n�=6Y�c�iY�3#�U �s�㐊�T�#�_٭��[J���ԯ��zV��b���}�d�"lB����bb�&>�s��$�:]���j�d�|G���r�� QO#����Rǲ9��%��x�4̸aqxK�=LH��d=���8�!X��k����	�WH�_�+�b�*�8�W���H�K�6��^. �Y�+�n�$�yE�q��`=��u�_��KF����G�B۴J�9���ҿr�_�o�*6����_^L�F�Y18&k���c��{j�ʹG���2�c�u��@�N߷L&!���ρA�s�63}
e��W��ZP ������"��0���k�op�*?؇ v� D�c%y�x���4L�k_�=�<����+�2CC�d�
�+%��w)k�
�{�gE�?������ӽ{��e4m3���@x��71����~L���A���Y0��QMt��}�vL�M����.�i��O���O6�鞙=������;�0f�h�Z2ꮌ�}O��.{妔k��Z'�r�j�l�*��'F�#X\��� ���u�+�-HLb	�E���Y��W���K=2QZI�($�>��f�w���˵����ÅLpM���w Gk���th�k^?���p��B�KZ���ѕ~��7�J��I�fH0�.���Mw�h��S3�5T�[���Wb�.)�nAYI�<}}K��&��Y��]��(ļItH���\0�,���g�ݒ�6V�ݙ9����Ġ'-�����k{�c+,L��++^�q���@-��50t�У�u��:��׺#��*�Q���GG>Q��ɥP@;��yT��n��\G�``�_oV&n��U..LCz[��.�E�>�(�l(}��|�n���>�\�������5s/�<<Ǒ�WQ��˳�P�K���'6�~b:�P�w����p�w(�zi�:#�گ�y�eI;x�/�]����K;�S&E�<������8	F]°Y~�Đ�e��\ UŖ�|����Y[.cŽ�')��.s�cZ���y#E��2����ݸ�Ҩ�p&Բ�M�h��"Þx+Ů�f�,:�^�m��s�V��hH��!Ί����g[��i�'_��P4A!H�ڼK��"�jf�8\P#�8a ݮ~t�2�-�b��2l/�B��<,.����^�ؖ(ʾ>�����۝�#�~��I�U݆�0�~���Q��ۯ����W�{��$(w뭖�Mkӝ�O��5�8���_E}U���J�)j�J������,���o ҸQ_��X�pD��;6��<��)j���O�d�Y�=��ۑ�#]v����xב��,��&���s��V�}���Ʃ��4O����;���`�4��rFL�q�������af8�ΠX(���L�4�4����|����s�ձ�!d��?ͥ��R�1	��fy�S�����+�Z�`�O���B^'�����A�e�&!�/�h�?�͟�T, �唜�Ƣ4K��ߵ�����FR���(j*�oɴ1�h�j����唵�?���p=9� ��id�R����TK�8�k��x���[��̿��IC�CL]cnU�g�}��PZe}�\w�|���Z���K6xe�8�&�VI毶�lر�t$�H����4�����rGU�I�x�? ��7��Xy�]�~���x^�c(��V�,�mOeg����'��޲�/]��l���2ױp�y�b��=ĳ��BG^+���5��̝;��I,Ly��џ}F2ڇ��w��Y8Wn/�.ǧ���a��!�Kp�� �MZ�B���-/�����὜�Aߴ	�XP�e.������&�?=���4��>�2�QA���"���&!UUfH��?��1����^A.P�J����[�X��e��j����o�n9�MG��>���^�Ǥ(�)��ڄ����"+�÷�<4]n�r�UQ�&�"�Nt`)ǏͥV�Òƴ�<#,��J�j4�%�`�C(
Z:���=����{��C�L��w��ת�]g;n�	�������F7Iu��.f��X�IY��:�����l�l��t��b��N��|z�cw�9"fE�z��~��=/+�K^z�AH�j����,�e��AY��i7xq�`_�!��+������y�i�ɰ9�2� ���$�,��Ι59VuW)��{��M��<MO����:�ʖ�N%�������|W��wd��b��|Z�b�MQ���8�8�~�����>KR��1�z�@��I|�X'�s'p����?�[9���?,Ni���<����MU���|�jnT|��b|ϸu1��D��4���v��������D���Aim�<I��E�﷬����U��.t�r�0�h�Xh���
s+?�W^�u����O-X��)��P�}���V��>�Ue�ϷP��(C2����B!�c;\ך�Yi�.u8������k���A�sT��2�a�Z�c�VZ1�r����g��nWz�9�Q2*��=�����{H�Y�����2��[�Na�m*�(h����G�Dͬ4J��_���Cpn^3���[沕0+�\L���F���V�Ck�7$�!)�E�#	�D�@�1���糢[��A��_@[f=�,�6e�w�@��{��[V�	��K��O}�R��C3��,��*�WJ�/P��5Ԉ���ሰ����� ��L����I����-��
��^Ƭ���8�ҫ���ˎ��SC"�WT�+=�?�d��G~����g}��[滯����ҬM��{���N��)��U�a3 ,����.�������/�����5�a���x��	j�aL�ћ�� %�发0�u�&U�����[��E�c$B�&B��f'}$��6y���Ķc��Y�:���ڨ�2��.��v��k�7��x*:��YqD�Ya�3�x?�o	�LO�c��0ay���XS/�MƤ1������}�Y�}$x7�ײ!h���_H�L��)�Z^�%G'�D�:t�Lk����%=�������\b
"�f߻��E�gl]�j�|-���mV~�M�E���9z�  �� ܲR����)�X����1z��>���ǋ���&2��s
��8���;d��sM��ؔ���PQ�Aѯ]u�-ѕ˨����%���X��~��.�_�1Z��yJm
}�Rv����[c���o���<�%r^���S����-��X=5�g���vi�@�qr�t�ҕ�cw9�	ܑ���%��@a$ۓ�u��aD)��#�D����ʴ��E=�
���y¢��"��
Op�?T E�,�,{����;E��)�6"za)U0�i���h*۫����0���)q�dA�3W��V�9^��P��.����4a�4y�ΖKsa�+C�j��ݿ��Q�U�-
N��m�ї��=ny�~�����p��[�,�!�~2�U��\����/�.}ck�+v��$�i�1~�`��/ĺc�d�L����-8�D�TjMs>8��L��e�>������Tt�?��3!�"�%B���2Op���l�\Z>fH*4[E�E@��Ԝ���G�os��I
�zF|;��
�����ot*�7����b�k����Ҍ���{�������+��n��� /_S�'��m*���-��Wv���A]$.�#{��j�Cx'��jd���=X�PX�͙H�Ў?�^�J�|A��!>�p�!��^��@f�,���e �F�Ғ��s~u�.*c- 1!ړ��9\3�M�81�E+�٧
o\�p���+���8�3��׎�mܸq-���cv_q���pG��Ӷ(-���Ad��&����D��V�,K��� �Tbڻ�H���^V��8�g�R���9I 	�j�%-�p�u`�6�h�b�!ZF�v��T�d����=,H�wA�L��x��~-u����Y61���`������BO~���N���@���I��ꉹSp6������)�+w��Ū����5۶�!���샏�I�	��
tU�M݋^�M��Ur����O��U�pΌ�?VW�Mg�u菾�Z���Ty�A��Y�L��
<{O��q8N^b3u�(��Mh�>�KfqK��u��:R^��m,~fV'`5�����Y��(Y+Xk��e�����Xu��Vv�ƀ�S�_�4���b�ʋ$�h�I�GX�w>'�J�]��I#R/������b�	�Z�F��
�'OJ+��������WjO��<�� �S
�f���^V�`C�K��@kR����	�{Aӆ��n#߹�
��xWs_0�|q���&�8\�Ʈ�l��C&�++��a��=�h{g�KtF��H��
 �u�aSo�<F'>�=�?ބt�E��!����JZ�]t��j2}a�<uY��B�z��c  l���K�t�2[ �B���W��C��$�	��Y�I�vs���D�a��4Y眽��ҥ����xz�Q�jC/��Z�?�mws���}�`�\���Sj)�������w��.j��Wڔv�r?�)��+w�|E�g��3sj�
�_��ظ%��#�wgٻ�܋\�?�ٷLW}V7���%�?z��Inup\kn�<@�Ɯ��c�O&@S�7qI��-eL0��'5Kv"�n@�D�⧡�g/��aW�">ڧ�J^J=����m�br�+蘰i-*������W$O��ԣ ��y���Z}�Z���kÀR;�%2w��ݐ��c��fڅ�[(=nC�O\��'���@\<�a���MB����|	!_��@h�����>�R��l��C�!ՠ�S����<H��lH�����|�.�^`�k�X�g)����7 Y����<'ƫQ���q�_����a��&��4L`L��{k7��	��/Y:n�&/�����ߣQ�5��Ժt�[ b�Ef�f+V?I��S��!T�������wFk�*��c�U1�T唛x�r*��Q�M�����B� ��a��#I��"�Ξ�̳Q"{�Who�k3�R j�U��	��������7��G8^i`w�$OZ��S^z_Ij	�?< )Z��6dA�bWl���2�à� ��]`i���Nv�pzL�ѳ�*����u]e��M���-��=�r�5N�Ht:�#����Z(���1a+��e�r�D�^�W��������2�4ӛ�g�8�XOs��_P*;ĺ7�ak�1\?˷�s�X�S�,�`��F�\}H(�S�y7���{����)%���*"/�sj�;"bg�b��D�r����w���e4��
h�tjg�
��yɦ��B�+zpmb6��މ�5dť8&�-}]*�mp���f�Q�D9vɑ9�C�m5��d�{�x�i�j�h�+'��-7[����7^�+�l�
Hn +��[�1����}�6�ف:��Nn��� oAt2{;|PU^�PPO��L�M��+��XF����B7|�]D%Q�T#�]¥�S�z�3~�v��tΡ��#���oz!���Q���i�UN��1�b*�4v$�Ey(�W(%�?�,���\��;Ez]	`��(�Qx�(w�vQ��d��^�-�ep2��mAlr}	�k���-(vj����{q��n�i��=H��_kڼ���zAOa��i����ϑC����#��2C�����mEp�0�Q���Cƙ�9K��Z�9/|ZL!�Ka��>Y������BV8��P?Z(���kg�����tO�Zn��M�A��.�y�k�/��[�wCE��M<��|WG�������/�[Ih�����{� �=5�U�i�wBEo�*/��h��f�*H��!�����w��9��	6��J�>�z|�&5o&M�)�ebMp�R[��A�s6���C���(À����<�M�xT䞴��g�m�rw�K0�&ݙ��D��՟^]y��0%���`�4	U
C�7I����� /�;P!�������c�C������G�n�CjX:� �̩�-�/)�_�6s�9ܯ޽f�U~��4k��ߪ��we�� �JPcߩA��
�z�������j��Jȑ�>�n�]5�����%ʋ�z��.\��$
{����^>~��-Ъ��#n�ط~�y`�����@�s(�<���^��y�L'��`)������y�3*�L��SIw�pQI�d��谆��Na�N��c�aU���	d#�����A*
!X|�dɣ���4i�'�����KSp�t�gI�K!�h4�u1�!|�M��珇���O}6������b�u��~�7���Y6��$��oZ�m�9����x���Z�=�������i�<����W��3Ї��|PE/�>��$��>c� ���Y>�	y�\���أ�#4w���&b�kƖr�v��w�/[�Aq����긷F;V4�*G�?j*���hD��0��b5�s�֨�I�f�'C�]�(��[Z}a�&ӯY��-m�)x��?�ʈ��"� 8�3�`�rt��ԟ/
�h��?)���7�^ ƀ�^�yyQfX�>���I��A0J�;�)W�gu�2G��O]��N���ߞ �úL?�N�ŭ�X��z״'�Eҽ0:�2��ݧ�"�h���{��OC�@��	ȳ��$�=���^'ھy�ﰀ�Nȯ2  &�i�f�+)[2Z���M0u���M��tM�ʻ�@��F ��\�y��4[�]�ds��:��f������|(��޴�%�J�3�����t���mjJ1��)U��˥g1����f����ԥ��b���QB��ɘ^Jr�e!X&k$*�sj���a�V왍�y�n��_��c�q�M�;؀n���S1|��/��P3| �����]����D8�L�M�\�:��� <���3���q�<T/"Yw�zR�G֜¦wr�AS�n^�#�����̑�.����Z@
��������ެ�W�W�"�pr�B�h!�>[��(�%#��d��#����,���{}H/Ҫ�:�
iځ�|�|�p!�W`�R���X���װ���&	� �z @f[�"�����J|wQ�)�z�*�f���=�w˷j���ex��R#S�>�B�nU�"��̗��&��(e�P���@5��n`7��D����ۯ��ܑP���J�M�=m�w<��;?H��"�g�t�k�C}�$W���E�qh�C7vEȷ�% V'�V!1��{�-gc@�fR�d��e��.�N8�L���b��4���D�ݑ7Q�\j<����9���5��_)y�eE�lbU�����֞7[�q���	�	:�,�O���K"H0��S�s̥��t�Ϧ�v����Z0�	Z-��kF8�z����[�j�L�c���׳j��B�^]��3+H膊���K ��xҊCl�� IN�^�%m3��ta慜]������{�h�X?�!�%n8�
0n�s�T"Gm�a�3�p��5>f<80��>!n����gtkMX��<E�5�Q"�N�4
i+"��E�C�����p�T���X��	�qD���m�)�<�'*<���UaF�� ��`4����Ϯ�dN����q����"B{|�2�6_K;�(�*0LI�	���7�T�
�P>Ln��xZ�����o�Qe@N���?h���_c�zK����Z���;�H~_}�ɪ�~HO���j»�7�{w�n��?kz�;�Tc�&
�i�\�Φ�_./N��9/ăp���|� �,�~���KqI��%2Ħ
�^�/��s�'獎�r���VIEg�t��Fn��F6V!җ�H�hk�F�P��(�E�k��rs+*Ur���<�t�.B��F�G����g�`�ٵq*`(+C����M��JJ�9nRr7�G0z&:�G(�Z���ԡ�����9Q�ei	dC" ���`��% <̟l��sM��qf�Ki������U|>�w�~��3~rv��]E��a���H�4�E��1)���(<�:;���vR�5��֎����v;��R�y���E�.KD���V�[�V�wM�q]�o���(�/9̬%}]�/r� @w�A?|��A�q�pt����4ZRK ��'����đq8Q7;�.��{`�lX��3SQ]�ZL��ֻ����Z�P��_Z�������>g���N�] W�D@8%q�k����%����q�e�2`�d���4�����l�H� _I.`��N�B�X!Z�xm�]p&�rG�k�t�H�aU�Ā���q�#��|�Elaץ�+c7��ܴ�)��*�|���>�VZ��\0V_�
�	4G/$Q6IP1��,�<��AH1\�4��dW��{�Z(�	q=�i1B��o�x�^4�U
XM9D���ҷ���۾���
�M�5�	X2#�l�~��Uɱ�<�AV�+<��(�l9%Қ���~>��ğ��.�K��At$[�Ê�X�_�O�xv�\�Y�F:b�L/��Y��/�c���Xl�V���?������#r;�:Z��;h6؝Zd�[�f�C��	D�bf�@GZU0ie���i�2F��*�!Bw�{�.��p	�T"߭���zma����R�����[��2K^<���,u�cU�c=gܫ����U~A%fQ��=X�t��:���f�6��-��q)ˎyI(�Mi1+H������/������8X��n_:�>L_��n�wJ}����
J����
~�Ʒ7nP�:-��3��&J�
����8p�I�k�Y�!�F������<�
�õ�<cWcg�������'��6�+���\�Q�Ò����E��b�J� ���-���Q���'��t	�8�+����uXT׃�����3�BN�u|P^:�ͯ\�0T�̽��d�C�w#P*��*�����=D�?im��� 8��Ӝ�%m�|��f�~�� 1=L��p�8�2q>����V�{܉P���&�Ml���j'J�;��f�O�,`�娝�&>�+��A9;���ĝ(���+z"N  [�W�ܢ�&�d���h֊	�#?H51:`@�����Q��m���D~Ow��aKb��+�@H�0=�����\V��m{�+H���*���g�r����|�B�4�eCn���k�{Hu��~FUG̾]�e�PT��G.�Y76��o��z�%��Ic�����Iޱ)Z�W��,ل$���̥�l�@XW��]L�ص>]�#�轗�L¥N��󡣔9�kd�a)Υ�P�"�G�s,��r�K�ީ��6V̻.��U�}2զ�-��Y��_z�����4T���'c��p)_�9��\�2W&>�����<�sX���l+ͦ���O��0xN�c�W���6�`�r3��Ƶmޙ:�K/�Dތ!ޭ�"D�.Ug��0Ҋɲ�ŰT��W&�AD[}L��~���u^ ����K���1]-����c)�G��H�T]��:H�+э&!9a�D���i*v����0h%E�⯢4,�L&����CNnPWK;E�TĚ�5u��N��������f�޸I�p��eWWMy�u��;���C�!y.��ȅ��=�(!f\�Ed0�~����'���.LX�x4���Z��s?ˎ���UBY~Vy}�C�c�R��6�P�+iv˚H5tA��z1�ŘL��a�����|�~����
��!y`X�2.��|�a ��`��К'���%;#��t'�=a]xQPK�:&����\�\O��p��E�5S�~�=�y(5tT�����3h�U�=[�e�b�r�����^��@�Ҕ��� ��P���7���[>�iz���!+x���%��˲C'N�e�	*Jq'�� 69�a��O��u-2��m-��[^����7�����SD8B�|�gg�A���j�?�"�,p��P��fړs/��;�rc?+6GD�@�$�.�� ^�/L&O.yE�8ߣ7�=�����ۇK�,��B�e����L}@��5l�|V0��CI��w,���[����U�s'8� BR.��j��Ġ��ƿ2� 3�q�������"T$�,͡��E`��N�-�dɲv&)r�4q(�ס�ȟ�w�G5/S�!�H`�Ƅb�ق����G̚�!�0�[`M��6�� k��|��U��6�
5C�h�n���l&"�}(M������jKcQ�oC��)�Mfw�K?�6��%}4]dj�����&�wX�������֯��v�z�����[�3d�Y�l�����P�>ҝO;O���,���rb��j�*���!Z�I'�4��*<�>�<��Yt�ȱ����#�խ��,�&�y`���)��?�BW3����i�Tm<�՝�Y��L�p";���7",]ϖ؉���h��2��l`j��r�'�Þ��]��/YO���}�����?�F}M��v���6���0]�E�m$��7�[��9���ǎ�!Ӕ�c�(4�Y8Ze�pn������t� Dxm�~e\�Ъ8=����sS��u�Z��B$M�12C��HR�hv�b&3g�Z��&|�t���P�2�o� ��s9ep��T����w�\��8�W�&YY�B���(�>�b9�>�;rc0�$!��`��H���shn_���y�E�T=�`��@�_�@��<Ky�r��*�xb�|Ԭ��m	Ҥ~,�JT���_�";{��w��ҟwc�=b�?d���������V�tЃ=�������t)1�t�u�]�9���-�~�nt�V�q\E�\�gľB{M��I������?��} n�%�q$ �����e��t�.gk�g���̝s_xȥ��خ�p�n�Tk���R�A�����Q���w	���Ĭ��A̶P;�ʫ�7���Y_�mM3wP����pJ�31��ɉ=�̋�����<b@��q��ë����?��`p�o����K�׷��^����B&Ui�@�ۣ4;r�Xa��Ft9�V��� �\Y����/�X�!yߛ�c=(#���5U�š�*��)�B�m�Ur3����yM-)S$ߒR�1H#dϪ�(�6�7V�W�����Wgj�}	�HG�̫徰~����ٙ{������r��B9Ʒ��#���z[b:�@#�įm��Q��j*��?��Q5E����c�+@��O���x@��{?	������p�`��}b݄]y�=��S�����I/?�����[�Mh�Sx���H�'S]-�9t��@���ukR��F(g���G�AG"�&r�ût=�.�b��%Y^hSAT[T1g��\<qM:�l
j�0��n6�2'&�,�g�D��(<6�.�v�YD;���[*�]�s�S���ۻ�!a�Q��W��9����n[^4x���,i�T6��G������?=��ܕ��~_����[�O������a�J��i�U�l�K��{��u�^0Db{�x�[C��O}:�A�1�$T��4|�����Y-6��ţ
��go�u�so?����2V�r��;96���2}گQ�K^�I&����r_�6)���Z�"��Ú����EW������G�N@P�3�*ہYX)�QP���ߗyY`~��1}�����:6;{Y>^v
�mM|!�J�"L�����c���X��J��w��M�o����Wwm��\8vVl��K�Mq�i�6ڃ�˂Hk�Q����E`�����W�J�I
�5!�$��3v�E�kX_~9w��0	���D�5�;��i\�'pIy�q����W����d����^
�����0P��C�K�&x��ײbW�eϥ�s�]��Цd3�=��K����\ (i�yn�hA�g0Ҡl��Bp� *�k׸jo>� w�m�
�����p��P����mb��p^�� ^��u�֍`t�	 { '�?N�x�S�������m7��@sk�TpȆ��q>�\��w"QG�d.�Lݰ$�O]�6�.bkd�{��w�p�������(����#��ݍ~E����	`1CV���B8�@i4gM�&H��N��JmE�S�!<$�S�-��,Px��}������wu"�B�:�����$%;DD�>0fUh2���
�Iу.���e�Cvǻ�}�(��g���n�, ���L�U���'	��C2�|��S#�,`�W�Ϩ)���-��s�/�R��@����@# "u�L�-e�:��ơdj��q�}��4g���ۘ(~Q�Bw��X� w�[^�m�
z����1�c�y+��@���l����K͔*���A�CfY�	�#�TX��C�
9Y��uU�/������K������ː����O����T}.�|���f�[�	w)V�h��*uiR��4�D*邀6��c"���7h�No�L����9|���\D��/��)MI�M뜘�cB@�,Ud�%yl�0�"R�M������N<F0g���W_\�fv���|�P6�@��˲6�^=���FK������_&�-R*/��&vk�a��,N5��W�acV����v��.@(�vmxc�K��
qĨ:Ұ����a��s�Z+������#-k�4�_TƗ�Y��#c93��Q%�ik Z���N��7�J-F~��p���
� Ѕ�|��'A*��X�dd�����I^+��(��K�����������
:��W �k J�Ňo�CD�>,�`ckDM/�D�Q�X������c��3{�f�����a��6$��-v��cu�N��Jv�+�����m�5�;�xm`&�c��W��C�H��l�X�t6��$G1b-� ?gʇ>�eU�դB��<L����HZO����?ݷ'���oqЌe��� |T��T睟�,�@3%g�h�)�_��8��j!����I�3p\��'��pG�N�h��1�'oN!�%A��������^9�ҤB�c<fpF��>��4.�E���Ԭ��{ɴ(��s>��$��`�o��rX�[W��z���t�[�c:Zf�,qU�ܚ��B^@=TX�@����ةS��~�HJI�2E�k���}hN0u�s�,�'y�;�ͺ�>�j-�A�r񣒰*-n�B����iKe���>�[L�D�ݖ�@���,ɕ��@F%u!ρ��D���$d�u޻��>ʪmGAz�6,ɱ͌9��_�W�O��ݲ��:VٳZ$!�e�-�"ʵ�6�i���G�$����m*ە��N�q���#X�;]�B�/m��3�)�E�l��"���ɽ���v4�����;��ȳ��M1�>���!T��GB�����:�;�V,�Լ�J���s�9�˗MsיC' �Bբ9�H�XL� �v��� V�V��<�^�>̗�C��xvǶ+��� ��*�&�8ک�o`���9W�67�Nێޢ�x�a������於��߰����ϓ/4𱆿��}����F�X���r���=�ʌ�4ᫎ��4L���������qÿ�>ڬ��V/�ǧg��#�=�$6��%B�;�9�ĥ��Д_��|��Z�%���WVE������2􍀄�?��-�h����)u�b?� ���:�eJ�����5"`�O�~���=��0�,����\kS���Y�t��V�mw2Z7?kx�_*��d�dܷ"Ђ#����Y�k_�sj,ծ��Q��1�4+�<��H��dt����I-#]Y�'������n��ȵ݇��;3��m�e�{ ���ܬʭ~�����B��m�pe"I�Z/�%�-�QG�aP�D�s��ᡫ�<dN|y2�j��E�(��'�x��C�d9PȚ5���*�5�8�א3��ϱ!!�V+K+ߥ��wl{�{�UN�d�Uj/��㊃���XE��3o?�.d>kf��	���$ZnU��Ǳ\��^ci�ݜ:����~r`��э��9^�!I�3�4����u�g������σ�B���UL�w(؊�W:��`��**e*P)K��4p���zό{�L�h19�������hUƃ� )X��if�v�h�r��BO"	�{Z�35�P��@�k��'��bD�H���g��2S�Μ�H����v��:��3l�V��îBq\_��@�����Np�����CO'%�b� �Ҭr�������$mS:�����*|��@�*�W�����d"v��rE�v�m?k���#B���neV�G��; �iP�L���sٯ^l�0�Gh�s��6�^����Ni'h�z��cq6�k߀��skK)Njֽ�[��� bqW�yݞ�F)iq7���*�D��.+}�w턳�y:��v�iy����s��v��D�2\[��i��X���c���h&\u����,��l�a�y��f~2#N�W)x���(�z� L��e׈���d��Y�	��%��%ZvSD[{ޘ����5�
���`��'䫗P�U
xwQ�z�w�G��+3�uи�aP\��M��ue��I!Q�������� �ɳj����C�]����D���d���?qY_��`�Xi?gc��Y���������T�n3�+TiKX;x��]i0��G���p�I�� �ܹhή��Jq�ȳ��wI�O��h�bP��Ai�^۶�s;M���K������dm��A����6�7c���T_�B�ʡ��^�C�iֹ>u���3B�*���h�ARc ���^g�����(��+�O�j!?���*��<)@P���R��BǬ�x�f�M����$!q;��I�L�!������Z��9B}�Ȩ%�u@8��H���\���Ȱ��4�ϊM}A>/�5���n�<�M���������Y�F�{������ `���)��W�K�Rh��NE����ɭ�OHK��D5�Zo�� �?�{���d{���e[��f�{y[���ݛ���е��0���%�N�C�u*LY9�A���ļ3�"o��l��!'w"���S
����i�jX��In-��dMV68!0#,e��^�l�$C��*��������-� ޴3Q�I	��gM��G&RL%�"k�VI��%�rjr�-Ҷ�q��)\����\"�"͗��/�+2�/�R�D��C\�cc'�7y�f>4���$��rD�d�vt�0��F��nrkA�/�i*��Y���m�;�$I=U���=�	[�]�ї���e�N�Ɉ�K�G�
(	oa�J�b'��H���̐��g���0�=Z�T�h�
�m�9k��b����x�Yb�6�8�ʎnM�A'�&���Q��/���RH�X=O(�1�?�7�?0�,��2�Oٓ��n������ k���{�[2�d%�2T�YʚV����뉔��<�C�۝Z�JC�O�X)��_�l�u��?H��_���.Iށ��J��y�*v�{�CFJ�Yr�ԅ�Z��]�e�󝟭E_>��)5	� k"|vd�IZ����ّ��m�u}����UO��rJ��A* -�;ه���tV��<rґ�MB�e��X��6���-�{0�z@ƱM��|��Ѥ���Ke�6L�^�Xd
��]��������A/���	��� g���ݤ�^
j��$A�Zԏ
��6��ny��6�r"�'6x��8����=~�ML�R�ڿ.#�o�����������z�D�q&8�G"A;1N�u�NQ;ϙU��A!G�~�,�]c���mS���h� &�*;J.v���I�U�N���:@e'"�����I<k���X+�>��WJ<�z�굋Ef��?������tW�Q:V7S��t�K����W�c�4���Q��)],A�d�W�Hd� ���f�����4�J���y U8�O���GƸ޹������e$�vV���J���L^����6k@�ܚXLNMhJO$��+���z(p:x܀ �G�b�"R�����n�n�~�W�Q���N|=�j>I"��2�6���X{aΈ�aul���IN~�<1�F��=�dwV9v�Q�b�&\�E8�syp�jtVEE�*�V�{�v���B�?�)���թ������o3��0=}�:LG�X����7�6땦�P,�b�W�(���M-��W]�!?h����4���)-�=�i���hځ�X����c������e� <)+�`@B�l VIE[���r����d!��y��'��Cα�2Mk{l�����?O٥�&�hT��B;XA��]�ĭ� m ᙝ/�'q+�]�e��``Ȱ�Lę�n�mS(;e c" ~�X3�+V0q�8Y$8�S`�͏>���>^3��+/��T!7K&Rk� ��蒹Bߡ����l(��:��OW�7W�}�J�`�G/k���؋��'�I�+ߵs���AbRi�܅V�C��`�^5bc��xt�<s!\�f���^19@S���!�t�Y�I2�,�s�A��em��h2�m3�E��=͞ ��z���$�nm<lO8���?�k(���?b�`�p��c��y�K�S�������?x��ԇ�u,,T"]�Ë����i,%&A�~l^&_?d���7��\כp���k\�S��@�˰���Į �I�05mz/�����9v*�_�J�>f�N�=��dh��S�����4�\Z;K,���Oq/s�'eLH�����Ex��<�1��jS����窉U���%p��}�����Co�o,p_�Ƌ�&���E6c����H=HJV��5m�e�We���������/ip/蝹��c��N<W�ﶋ��=�9��I:i�+� �V@���#tH#�Ms|G��^w��+��*�WRT3���������t8F(�r�k!\�
H��u���F�/=���V{2y���W�u� �FM_J���|G�� �=g�ʓ��$<F]�Ǒ$�6�/���ߔ����	�c܍ ��*ߠ�>�&,��2\�Nn��s�`���4]eT�J��?ymB:%������Ċ�Z�)�}�Ij�Bx��.af�V�{T��8�@��orK��X����Dg<NF�������F��b�T,����Ǉ�Bu�#G&��iimA)��h�#ۜ��䒢���3�<�H���*`�&+��p6}j�f�L��i��~#��	�����%�CՁ	�x����#�����
A�#MST�y�����L�n)Y�
��^�W��$�Y��o�4���Q+��S���C�	b�����q�P�|B�����=�Em��P�6\Zϵ�^����{�OZ�`'��t\�J��ԑ�!X�^�F�e�A �f�O�i��^��g����K%Jj���y��x�c�6��B�����I�C�IGM늻^�E��l�g5���r�4Ҿـ����(8.MF�cj�B,e������9>�_M`�����V�5�׿s�BC!�m�$ƃ��M�mZ�cE:@�c��$�{�5���J?
���E�kC�r�yU�Gr8��O��$���\�j�,���z�"5̾�hZ���%�����O:��m/s�Z#w:3�.X۫����,>��iAy�� ��l�d^S��m�[��΀�Gy<��n�I���H�������7�$��U$TB�-�3��}%��8:�������+9x[�!�o6��5��Ud�����Mw�ijP!9W0E���:�|c���7�d�� �����Bs\���C6���QB�ln�aUTR���$���lC��:�"��RXb)�xl�+_���L�l<#E�G��9��/��5��E8jSP��!��Qt���:��m/P���q��52_���ŝW����k���)�d�zk�&c����צN��f���|��r�9xJ]��.�S㝖�|�<~�i8B �㻪8���>F�N���nZ�6a�2:��x>�}�{��G&8
���W��V��鑔�۱p���7�Hr.����@k�i�럭�R;���L�P��6@cb��9�ja���1J�0�H����u���ʭG���HY)���?Y�����U�$F�B���z�Bgv;NC�z�:*1��K�`��g�+���ܧ�%G�l$��E
�[ U�F~y$!���Rv0�yBeq���`��*XF�A����0J1���|��jqC�����g7�#���h��2�)���q�#��D�OH�܄�/�P�����S���x�z�� /:af�t�7p����zwR�>�yɀ�WD%��r2�ض2"�A�X�2������B���C#���#D�m���R��e^��LKI��@
&�QP����m7"���ze�W������+�I i� �yI�mᒔf�т-��Ɋ/��_q�M��)�q?}��#!����.�P6�	+�\'��*�@���KxCI����l���즘V�`صAڂ
'(�0ڵ"|���ME�N4JA!8��td�}��aۦ-�O�h��H�N\��߱�H1��>e�x�07�s;��&�Ċ��}�N�I���nӶ�'.G~h�o���_W������'���e��&� ��f��)?�t��a�!�0�`c@���H]���#��\,���$�]�����!�b�qW
L�v�.��P}�|��Ġ��C�C}�ᦀ?5��FTC��@������`R���<�`���aM'I���ꊜv�N�6r'ћb�M�w�L�9��Ԑ?�V# ���������_�	AS�֫��Ct�.�ŵ�M�+�Y��M�)�K$9�m�d��C�%O[�?C������¾YMC�%e�(���(i�ZC��_W_��moAkVy����j�x쉻Ky�W<8��՗D��KJ�1���=I1T� �z���o�]gɴE��ת�"]M*([���s\E� ĺ9l
���r���KO}I`���r߽[�$��6v:ٝ��"iE�����G�H�u��il�`�WMi��?q����Q�.�o���$ɾoMj��#��~�r#fqW���nnE�;C�(ukiS�����V�lvf"�bӥ�6m'��Y�p�Tk�w�v׋\�!U>��x�Œ��?�Jީ"�Q��x��6A.�g����E~���c���j$L�+�Qs�B�Ɓ����9��4��b���K���%SV�ڡ�=慚vqc�s���
�B|�/N""( m�x��U�<�����m�*��?7Z����Jf�b7Xf��\VbA���%C��������by�;:��H�6���̜chY1��������D�5O�]U�y\�&PT�N��t��̒��x���؁}pO�ky��'��^����?�*5��UyC�\�p��Y�Je���?=f�K�vq��!�J9�J�N���%k�E�F��,~�.�7]�@E�c4��.���	0Z���DE3қ�p;[��̰@��e@Y��5Ж���4H���!^�D���2}�&��si�C��A"[l^2߽
�KM>�
�0�K���3�ʏL<*�mP��þ��9"�V��9!>���Xw�l���㽗�n,����8"�75�~�b`m����ɛ�g����4c6��r&��eI��z~������m���g������wv�W��޷!w�Ы�#"�aLY��zwS��j$�}ս��	r�K�ak�u�2��+H\΋�;"m�i�Y���ޱ���?Q\*�+���Ȯu�0���I��j�r�񂧨�K���=7�Chugz�����.��l�2)&�	ǥs��f�^��W?�U�Ҽ	;��o�4�}��e�Y��*]y�Ua:��,m�@��G�v�~��
���S2Xj,Dk���}�<�$��	�bf��C�ȱ_,qĪ�l\�w՚���`��/C� �V��N.|9D��.�� ���3��VNF�!�z�^�B`Vf��vT):f���s��:�q�I]@y�"��+ȁ�!�T��.�&!���1^"�H`#�Ȭ�S��p~�E.=gU�L���T�Ӷ����-�F������I���,�����%������[$W�ۙ�,��z(���P��J1xJ5>g�9:��T�\�i�啺7�?�
!��w����S���\��{Mr��M�|Z�����*�\������ӥ��J�|*
SO&*��f�bَ{7L�����g��'�O7�C�\0" �{���^�r��pI���?�鐇�N��j��8p9��ӛN���g���ؗ&tG�f	�R;=��%����n;���*�� �Y�i$�,3怶��s�(!jJ�}yz{F��0�9�|�C�O�'���*�;����(㕚9�;��
�nB�[��Dۥ��NF����M��IC/=���h�@�zM�G���l�P�m�u3pD��[.>:�a��i4�v[�J�ZC��vw���;	o|Q�-�YE�m����V>��MαX��Yp�����#)�-1���Es���pv>��[B���y���@��^S��S��m�
�*�\��jB��9�9�9����2&pgwՃ�m��8��1
��۽���S�!��%���:\@�,���|9V"eπ����������4�1���=�~���K����Խ���kht�S���}�sbyO�H�w���}B�@����;w� ��@"o�!t�YM����	z��ݲ�	��e�N�lV� �J�!��I�����&�Rग़�^/ϲ j;U1��ʹ�7��*�UƢ�g,�����󠠝�Cs�BQ�0�h�����:�@"�X�N���U?��ܒF͹�o�$�:|�12ڇT$��,z#�#D��(�u�\���y�%�s�*�[EO�~`�J�_Of,�<��S�_����f&�\�A��`��ܖ�oS��w��z��RF�b̈́aU�8���K���v�QkA.k4_��|L�ݓ���ºU8��E�1�5��Hńt���H�!D�Uh�5hd�?�e���L#�.�"��U���j�(��qG�*'��]�t�����I����=����>�cH�K��Xڅ� ��#�@�۪/k~ �9�fd�=>P6�+�G�`��m ���xd-�(��ڤ�#��;k�6�<��5,~��	c8�H�
�y�|F]�?]ԙKdǄa����M����w* �;��࠿u���!�m
�i'k���M��W��O���W6�b5kCܥKB	s���ߔ+���[��q���E��l��=��+�)8�I�L�������{|��DN :�G�zץ�,�O����%�D�2���qn��4���o]�t�:� O"�S�'�2�n�0����c�ǜ�$�&��؈t�M�kl4��M�<8��E������.��g|^��Hoբ�ʖ�٨�����	��u, �}[	7�@P��Z�I;u)4������X}=<�>r82_�1:S���<z
h�iR� Ғ�ql��Ӈ�����E�GKpti㇚�fwS$�/�}������H��
�6E����	�.ӧ6����7GP�t���C��iz�
\� ������P�2����-
� �-�Ġ.�����S6u4u7�,�8�:אWh�B֧O�#�*�PB�� ���oӏH��5����C{a�cj�3�6 �b��oа�e��IȈ!�~@�)�n��&��n
A�M ����C�����u;
��>�`�N��Ph3Q�˱�M㲂���`���/��A���u�DJ�v[�/�s4д)j�jl�I��
zS�� x��\(" �"���2�*���Q�U{��k��h5��n�֬3�F����f�����=�_����/���.c�t9B��V\��ش�������6I��`/�:E��G
^
K]O+�9������1�>�婟� j��}QoFkq)�B�OT�p@z��ray�+��%�)�!������~F^�F�܈�4�̀9x���U�QYɩ��pΈ�fb��=l��^��LYXI���u�Z2�%uU�d!Ŷg��}Al^d[v"�a� �u�sWd� �=0��}\���sZqnV�J��_`�"OF����j^V��������ۍ��B�!Ƌ,���Y]�_�&�!7}A�Y�����c �,��Ji�$��g�S���K�zy)�S�{���vR6*������7���x��̂�&�H���̿LP�0HA����Uk��'t��4��V��Z�ړ�8�ˉ�^�%'a����#���w�a�Ri/Eu����/NG�u�i��$C�&ͦ-B0"�V�-�f�C��m������|�8桂�xm��n��1���#��x(ʉ*Jl1�Ǣ�ܶI�*���ahv�S�&\$��]J�I! eFx�(��~j�R<�]�wyC]4��+���<7���K��Q��6h2J
a��!��<�g�+��&	�3�d��k2$U��ʓ�_�Cj�C�Y�aT+M�V[�=��Eߛ����BV��T�AŹ�X_*�|�tiR�}Q�jyh�O"����{��y��p�Y|q&vX�SMӳ�%嶕^�{a��c��O���z�U�Ѣ[Y����̡N�xf���:;��Zi5Z7,ԆH�*�GR8��n?��&���rM�o���FGb�;��寈^�A�h�q�N8�֐�p��2U��k��d���h�[d}1W�T�T8|sd���"�r�Dy�n����UG�~��P����O�qs��bWory�#>+t�$w&4������A�c|AIW���Υ�S5�j*F6��l���x����C��U��XГJY� ߓ��@1���9Y��A���U5�����*�o�H��#�ihl��T9c��ۅ�}�տ�s*T|�gt��H�`"���;�8��y{}/B� ��~jr�O {�UjG6�2�՚"��O8EX&߼9�]��z���f�43��%"�ʕ��}%�R�T3�@܆*q�fr�{X�8h�D�xnfm� }BP���8�ճ��e�H��G���6�����B��������w�d�ڶn@��|��
oA�|b����M(�|�+�goG!f�!32'{Gc�2�=Y�w7ߏ�D��ZWI8� �19�k�QV�7E ԴR�kC#�,9Q��b�"V���}�&�fR��~�IO���C��2�=�{����JO,]�k�C��ȯ�d�̈\��2�ԡd�/������c��#�����_>�-^(>l�؋��P~�3�ͽg�(�e֔���D�ٿ�^,Z`
����s��+�5�y�]��+�9�����
�w-^�v(N�b�,��o����IA�H�����U����:�`Ʋ��$�b̐1�F������Ί&��vM��5*��w����	�s�V�:J;��@fM��;�\�%:��c�nwZƟQ���� @����� udE��?;�c_?v��h�LX�s�jn�om�ܤ=��浸��'�:�>v�U�)8m�Y��˰�O�K��Ҩ�L
�d��E��2ܵ�|HYn����x���$_�է6WLq����Ԕ簺�B� �O$ČJ�Z�w��ir�[S�<5hz�_�?���w���^QXh�1�Z���8�3��v�?E�d}�]�����!�n�sz�@����:�3R�V��F=\k:��ޗA�E��yT@�O!�	c��!r�w��%��2.�9�H@e�I�5R;���B�[����ܒ�=!�P��'�5��JW�Q�
�֊�|��4�YЃ3����q�O����s2y��>��i�ܺ�f��Ԓ�>]=�S5��?+�hb�kI�����8�Ef��P���^nR���;�2�#��(�ܻ���m�~\��8B�c����7z%m�B̎���Y
�M��@�o�Q�I gd�������ݭQb�s/i�)yN����p����Yv����s%��W���l�u�������\]�1dP��mJ߉A�)�����zg���΢<E��1�־����Z9Ԍ}�A���7*^�����cH�I���������{�0ԏ%gE��Z�b����Yn���������A�;�V3W���ۣeكo���D�d�=n(Ur�ɯp�7��`�I��7wxP��ٰ&�'@�������Qj&��q(�!�� �ތ�j��1&������6�v��c����E:�[���~Aɴ��%�<������w�dr�gN��/��\|��s���`���h	���taՂ�a�q�mv�wH���m�R���(��{���}������}��|y��I�#��=�E���[��-5÷�V1C;���w�a��]m�#< ?�[���G/UZ"����iX́�������F؇n���"<����ZHx��7�K,�d��)b/�7�����uY%�`3d���)_����?ޮ<��#:m�u�B�IV����s߹ƙE.�<p���ړ�����ĸ;1Ig�� ������݆5��X%���i1��p@�Q��[�⌸D����S8�D�Kyq�e?�ؤ�7����2�MRE���ά�I�4�K0�D�B���$sH��[����Κ�H�ӠcrkE:||�y���X�gF�}�$p��ܾ3!Z����K��ݑ��K7��FI�0��
�j�4���ٓO?�&e��'��D	�ˋO�n�������;&@*,c2��LdW�GU���%v�=״���
J�rj�S�g\½���������7c�P����)��{�(d�2@~���ғ�Q�� �Lk�;�g언�cW%��-�A
,�l��F��}�@zfkbIû�d�vr�3(��Qc���7sE��23Cc��O.yŹ��=I��`NmK������{�֪�o�к�G��� ������Y���O�5�n�9Rn>�A��vmrzk�fl>E^~}"�%NH���|%��o��-O��/2U�3�7i���p=r�.��J��e�sR1]��f�Ė�_��Ғ����X�;�'N��oߪ��+^�5������J����4��O��J]ؼ�:A���@'έ4=>�$����� �=�1i�Q��b��m)0���)]���'xJ���Azz�H~�����{Er���?�cc��^��-x+����q��Ǘ���K"9l
@s.
@�
��3��<ɸ�Y+7�`�{+m�Ou&�=ٚ�l�R0�b�>x6s�������Df����p�f,K���nH��N[9��������m���S��<��|�h��W㇢[u��,�E��]o�;��MK���@��th����[��%�a�����T�]���~sFQcʌ��Jx�@zPP*�ɏ覓�qG��ƅo�����������o�m��?s8T} ��
p�g �����W��{���U�
��Yw��^Kޜ�����ݛ�y��W�q!���/T��]��={J�JA�|F�q~m:=��ht�U㇋� �U�	5��~)�S«,��;旫��I�t*e����َ��&�2���Jg8(RG�^���������)/�Z�q�2��1,KLʬ���d�|�A�4F=�'���4@Lf �z
�l����o��~Y�O����\e[Rd fô"�|Z��hKM�����9T:��b���� xo8�Mt�&}y2��!U1�7E�W��M�t(R��{���CM�/�V��űR�r��t�8� cnp����i��Zf&-��
��Dh����Z݈뵇�.ˋ0+Lq*[�<~�����f�˘��
gTلW�a ��b� ������Ge�pD����W"� �+�&'����qsxrF�W�P:oyـ����Z��y6`�.�CF�o��3��ύ��ވZ�8��]pva�ro��	
y$����e�E���I���I�^|��z���0G����^������~d�(�*y�>���<��V�V�#���4+b�*;6�����|��/�L���D���o�j��Z3V�a!�u��"��3��*O�U��9���t�nk��+��x��C�����h4�}�ɬ�z��� I,0�U:���فpںlG��$-���+�Í>���&8>[��aG�ŗ�c!�p�sN����u#U�?ד�3��}f���z�`�ά����Sۂ�����n&<�qY6E��܉ 2�-�|�D���O�Kk'гڐ5]��Y�zk�e/�^��P Zd�g����szb�
n�.��{ ��'po �,]ݠl������2>~�Zz��=h+�Iނ������S���,�	�us.p��:��$V 4�4ю���kҴߋBwƅ23H�܌�]v�s4'��뺰�ǘ�����D��
Eh^�̶M��޵�����e�%�'wJ����疘�6j�m��t/�r�%׾�w�F�D�A�Μ��TWb3��e�?6LF��#��hD��P�*�M�˖��>���#�^pG�S�, ]~l����M{!ڝT(lx��)��0,�`(N�������]^fD���|������{Nu�����F�ʌTG�����z� ���[��`�"�1P�PJS����CV���C�Vo!�5��f��
���r��҂��_۱���]+����D�X8����q~y+��ߕ[�8#Ό��[��9�YCe�6w�M ]�抷���墋P\ߗsg_ɍmf��V�k����C�NX/*?� �.��8�|z���'��[��Bqe#`��Ѥb�5H�|�kZ��8�z.��$�¦C.B�c�i>)ȊJ��<�}X�w�4#��1�b����t��G7�C�V�]cI��s�p�"h�[��
9�|�NRLA��Ց=�@�o�Gz�5���#=~�:�H�����X�;߮�er�[�)9j���xm�$ݦ|Z��3��~�vŔ�19���ɶ���5r=���h�O��W��?��:CAi:׌<BF�жZ�|�*[R\��d��Mb��;s܃ҤQ��xy���!�tB�F|C�l�������}%��������ghA�����X_t�I�k~�'$[�k]� ���#��������m������u"��e ��Y�w=|����{%��M��<P�T�a��F�%t���E���|,UG[$�?��I	���	%���?W$�Đ�t�Ԋ$"�]��o���®�A&01TIp�#P���]�yb&�Q��I���L��O�2�X�����w+?ѓ>�x'���f�h;�P�F
l��E���B?�
??��㓫��Q��e��t�I`X��'ƨ�C����4�	]���_LYvH���0|��L������� �Klyps������ͽ�+�y��<�_pg ~#AW��B/:޽�>��#[њ)���hN��ev����l�kɊ|��Dh�u���*`��̉wz�����Z�F���t2�۞�+艸��d��9�7K(�G����@�;}d������X�R7�M:!��.�!�$�6Xܤ9̈́X����h��B��0N@����~a�zNDo��@'�iss�Q�)L�]ײ�\ٟ�^Л#w�.|xs�~�$	*�7d��Ë]h�<��zɣ7��@�a��bho�)Y�7q�;ж�x�����Gv5\K�G����J#J,��SS�57������sD��N�1'ojN�f.-�p���G����ZB�b���y�Vr��b��j��A��f��/>i�6E{B�錻��4n�ʷ��d�f�ᡤyۻZ]Fj�?Ϻ�Q�x�F��R�ZQ<����bҽ�Κ3�ӡ��(�
Y/*�}PL}_�!�������Ά����Rak�"Je������[K[`��f
�B�Y��9�b]
��(
5 _����F�L�{qOrP����R�4�*��ݜi�Cɡ	�PB��y ��*���r�&?���Z�@�[�� RuP��*̢�\s⦩��ܑ�[q"��omc
Os�r9�2x*D JrCs��f�w1�L,�<5�0��N���%�H�j D��ݨ�;%V#P�g\���О�~`0>��u���c���,0g���M��o��qm2�э�=o\��E�:h?�%�<�HA(�~���5,��#��tN�&�$@���̲(��|�iaX�ۜ��Dߊ����R�\��'W���"��7==�!2Eϊ�&1���Q��ؼS�o��o�ɩi% �9]cb�-�E�]�5���(قx2E�`{?���b1T�9�x�)vT�&8<`K��Z��Xz��u��7��0&7F�Bʦ�^�k�K�$ȫ���9j����i��e����\�9� ��C�L+�3dH��t��ߒ���#�=A�Z�n	 g)ƞǴp�h�ՏJUgo�FU6��doY���"�e<q|O���AAB��/R͂������^����:���y�v����>���޾�{�d�=��xS"w��G2-j�	�ʨ��PY)��Ҽz���t1��k:ק�=� �O�Pgb0����+�rv�9ێآ\ʭ������r����]��.|r���*��S	�S��9�N�0Y(�_�*�0.,��@�N#B��8����0�r�ʅ�Z����&g&��0&�p�,�X?	�������U����;G��
������Ql��ئS2;n?f�F��QS�Tr&�4�_>x�Y�ΆM:a��=h�����; D��"V�7Y/�7�@J�L�E�=5_B8�
��K���\��}D$���*1��z�$�������Ɣ����MT��-e����j�4���/�����=OG	<80gЋ�.	c�����M�`���+�O.wA4V��QR�= ���5�c��f�t[��4�O��[7M�^��Kula��X ����<��L��L��,an�K@�i���YF/�B�%���v����>���7�d?����MvҐ�D�G��B"$l���$W�R#�� 0��8�؟�`v�8 ]�6|ʟ��<?4�Y�{�9��S*v���2{	�F�h^��Ā%��F����==&�m*�'��l^�fks�m��^���ǻ3��-�����g3�5'�Vڶ��_���zI�R(xM��}���P����Õj	��[��ې0�������S�lFw��Tp�|���_���A@wJ_!x���}δ��Ęt6�,���Ys�o�O���}���s�j��~/���\3#Wk��
��[��{���	t��R5�w5,c�"WBy�^M���4�/�k�Y�~����op�В�>'��������V���%���fb�'��	�q�� }�+[��f茊�S��I�]�N�5�&�N��X�yD������������p��bHӤq�q.´�@��sWg�&�8�S@\� �������ru��D�7E�}0I��b(pE.?�zc�9uomZ|��_��{!5)j��.��z�$�"n1?�jr�!�p���H��~�pp��������sX��e�b�S�Y �z|)��bj�8~)ا��1ݥ	�L�H�{�E�9-v%��ϫ]��fC:�R|7Wp43J�p��N�.�M*����
�-r^k6�Ȟ�pcH({�fJo�"�$�Za/63���jo#�{\x�,��L'�=��׮���1mG�����I���4O��WR��tho"������5A�Rv��|�8Fp:��1��X�/P��O�P2 �����ʆ���=�Ld���,yۃ�]�/U��{v�_5�M���G*L �򫣈��DK��n���,�&E�To��Zl���s��n4�#l���@�J5|��^�(�oD� ݓ0�w*��Bao��Y�E�V�+���?�����g�5�˨��w��s��tJБI�b�1�/��	7�Xe�-D%�(��U�8��Z��ᨗ�M`h����s�(��L�KA@��h�[&������'d�KP���5��j|u�%�Y����2�uKꐀ4[6�e��NEP
�3��DO���Zn��b���.�45���3<��Uuw�����/��s�^�b��%�+�&����\LF8&Ũ�$c=�����������f��9��/Fy����f9\I��s��SϬ@�j��kP&>�V���\x��r=�>6;�+]��'nX7�УjKB�n��Ot��V�2n�Kd=����(u\��ݖ���\=����n�Я-@PN�Ϝ�.�V��Ѫ0�.�ϲ�Ԅ�gr���ΰ��!ܐ�f>Ι��L3�_V�Gc_�h�;��z�g���p�-cU=�\�h��8(�M��5�d�3%L���ː�N��`�Ro��Զ���rq��{#�HZ�`��w�M#ӎ�W?���s��Ҿt�M~��Q��VMv$*%�P���-��M(�t�.)��ڄN�t�Hk�7��C�%&�+�Cs�k��{g�G��=dVUzҴL#9wԟ/����9o����xɷϤY�����L���}���%t�L����w����W�7��\.���E�z�\����y'S�g40�>A�P��CP)^N-%ͮ~���_6|��d�g�	����C�j�P�:x�lL�Ji`=o�p��'�����-d��fk���d��ev�T�����Z���b��۾�0QL���q7��L����l��<��.���o�7� p�t)~����r4���J b,"�� �'L�-�:��o�QJ@��^G1����y���-����LeJ��v��]^�H�����J�Gțs��0��Qm��u��p�X�{�P�d9��bb�m�����P�m����l7�F-	�sr�<�����7d������*����!�)H�1�=��<�5��ҕG#�V�~]�c�����i�i�;g ]�����o�n7�MH�ż&���M����/�H��mDNz)b�s���d���۸��wmeZ�������Cy�,�_Z9՟g�d�'�~d�D�i�~�؇�v�Q�A�Wx��`Gw�� ���^~�-����n�9%m��-�|��#��5����Μa��_�Kz �+?qm���޷�Tdtܧ�iQ�S��؆VʭkF~��}�I ]!f<�W�L�����\��޿�e���v>	�1^��\	��ܸ����u~h����E�tVdl�'p��-�����Z쀳���L���S����M���F;A���� Z.��"�1�X^����������ٗ 8��[~[<r�k���N���ųõS'\{��M��8��������Y$>�5
5R4-Z�vfz���q|T�w�	�?�Ёuw�:b-'La���
�tݏ0ˆ���a��m�����G �gV���n6��4����V�I`m�p����0�� ��{ȕ���C��H���қC��n���ˀ�';n1���r��Vv�)P&�8t����c`���.	�c����4&�ȟ�J��d�@�,��%=�z��r�	L� \�oM���=�`�I���8\�8/a����*�g�}~*��Q(�(�r[Zy(h�$�oǈ:�N��#�!����J���jSO,��\cGl�������@�(�"���E{*�4�^p�)Ҥ�cc=m��.���U�l������Q'<W�.�$��V	��.f_����%9Ӄ⻨3�	�;��Iz\g�Q���>a�!��)P_�y,z<��|6�/�/CV8�.�\�"fS��F\�<Wơ��w���Ғ���1R`�*�"�@xT���R�s:t��~_H�IG��3a�j�\��{��a;P���z��d�_�%k���N�����������"^�/�Gݥ̴��Fg��j��+-�ԌFz�{��Z.���'��׆�������\�d�
�_�2�?w(�?�D�VN��"�52#߮``��q��I�ߔg�d��̮�E'Ը�U�$�gR� ��d��,��lכj��$�Li��������_������cBE��U��og-�h��Bp�0M"PJx��5�oK�qgW�JB��
Ś�>~$��zh�\Ί�Y5Ň�AWr��l��MC�8��(�-*uw��J�]%(m}��>e�Om��y������JQH�᠜I�э0�y��>��~2��a����k��D��� � ��R`N,�Si�1��7�j�Й
�ȭުӯy�*��!�V~x�,�8ptZ��+�����~_Z�4[��3��j~3a �:�cc<[���+��,-C��zڻ�/M��C0^7�_XfY�J�����\Ԧ��O�d3���:2m�U�J-|p༦w|O��Z���uUrNq襟�LWoZ)��rH�5��E}T��#�b�D	�M�i�)�� !�\o���<|����n]���_Y�����]~Rj�G�A������E�i{ѭV�N�o��z~a�����Z���r|�#������E�����K��K��T�<9��B�0�N�^�$pߨe��L�Z�os��a�kRt`%����'�U,G3�ԕ���mr����Odf%��YW�_���L���u ��fi
EܺJ����Ղ_s�컏��-|&���o;�>#`A�͟��^M뿗Zuն�����X�(UE@�ndv{���sbb�4��w���>e���z��f3Znw��#$��xߒ"�񾊥��}sܻ���U��_ʵ���R��Je��6E�%�~
 o�t(J}tb�)���p�`$|����M_L�.��N���ɝ=��˰����9��l��8u�*��=�G�s��-ҴW7;���gC���~�S0�oI� �fbFKZú{3�AI6�pء�h>o"�h�Ə֫}��n!<3+�]�002���=�]%��$.��s��6�N��@��K�s��Ф��g�{e	���\�s<~X�.��t+u%�y*n��qi�i�|��p@���~	X�Z�{zi���H����ow.S4�)��/a�{߯lrGp��.��<k�L.��M����H��Z� �
���_��,h�2����Ӈ������+�[) ?�>�3x�:}q~CiRXI�E#�H~	u3OM�y�5��Ga� ��)$�4���՜˫�	���Ûw���W�E���D���S��陒����aN_�=�Ri�W:�40VX03��W�U�[C�<^W���7����J��|+|�d�)|y����*O7���������7������*�ϠnwW���p����D�������e?�)}�Ye�ж>^v�2;S�U�A�d.�vrAn%G�m�"�$����]�x"��W�<*�8�E��8aWN��5bd@$]�*h����n��Q�%�P�s�}�����cb:� ��Y�k���X�z]��}�D���ݹN�9#R[���L k���^0�4S�|�ė���o,��&�\�Cg�;HL�m���0J�<>R���T�NH����lE��M�Q2��O�����<�n��|��e<Er򊷏YΑIKK6s6��a9�����5���/�u�	�#+.[c<*�����/��9��X��f�u[x��0x���y(n��1��Ӣ;@h��q���@N���������<����4�ݼ.�!=qȖ���ޮ�)��E������}	����I��r9����'��ӤMn-�k��y���)[,᱈y5�a��ݾ�ߒVװ�:U�n 9�F�$p�oW$GZ�����g{�� ����R7m�6���$���A]����뼎V��b� {~y��Ѷ|��ɶ"��BO੧m��Th��U�
c]k�h7N�Gy����y������o-x9K�6CP4֋�����R�\��
�?�����fb�Q� 
g�-2���+�۹���N����w3;�7b�DH)�U�qpհJEe�D�4�1>�8�'�",����2�)u%E<8�)���=	��^��j�qR�)�񼅳�7�����>Cdgn��n>8�����s@k�:r0{��/�Q�	f�B�B^9�T��o-�Q����>�tg����©�9�	����0QL�v����	{�������������m�z�uFBJ�˯~��ϕ�]�0���>W���Ϩh��#�K6�I�Tg^�7o�fF�����B�����ϱ��S"��I�	 �|w���:��߀��BV߄��T�*H�N� �	�ǫ�qWSf/���I�#��˸��h��H��8�8�\,� ��d��/؅�6֖�����FrM��h�t��iN���_�+��13#�cL�1A�+d���uୂ?��j�w�Nm�����"o5����2�|FI��Z��_�Ix���R\eT�#��\#D�����$1�A�������w7���kB�j��G1�2�C.7�cXf�*��47��ş�
Z}Q��:C��^*7��@m���<1ZՄ�S9+!N��S�q���(��9Z�3�GZ!{@7">G���m�{��%��iY)��T��M�(�/Xn�z���{��A��M����=�,��
 #���l7F� �,Ӭӵ9�t��K�HKmvX����pXBk����-�K%���m1N��,�B(���,��t~�:�vQ��z�������c
8F�
�gPƏB$.ljo_с�R4�ؽ"�=��L��-�{B��퇤g2+ӂ��q[����o<D���"Y�GjB?&�x�Uo���L�Xg+[��kM�]ZJ�A�����} �m�u�S�.TJ��b:���R���}�F.�Bb�Yȳ������n���ue��p��_���`�0�ì��a��(S7\m���K�q�0��L���2É�򴭓ki#E��K
�Ԉ�p�՜#�zc:]��^Q�I�w?�K4�+� �)����C��n��u6,��\�ǁ�(�{:�סe�ߌ ��ʸ�(�|�* ������&����K����ޗ����d���r���������)���0"Zs��҄���9KQ�
��<���u�k��d�>ۓB:o��L��D�j��_L���C�Td��w[ n��;�?�:U���y�.�-O\���t�FĞ�*��
�,Ζ�MGO�ؙl��Y��ֵ�#�F9'l����v�)�g���{��/����fF�ރM��g9�2�-��qڄ�IWn��?���P�kx�t�,�y�����(�Io��ŕ� |��6�U��!�I�_9�#��/��/��׈����z��Mҙ����I�~~���03�;C:K��	��]��w��K�;����&:�ҏc 3��5'���Od�+��z~�&�R��8�e�J����K��g$�/�׌1Rj�l��%8؋n+$+����I,���L�eüm���{�{�"8�v|�;���"�ik�i��4��*H�^3ą�����
�t�AH�CgJB�4�ͣ~oe/�� z'��r v�*ޅC�/>�lyW"$����U�8�5lP ��+��ÿ���X�!	Q�<�$u-Q���J)�\��-ft.m���Ƚ�8Ｗ0�0$��V[���Ja�U4}�6̖�껱�`��ӫ�@5ߝ���8CH��>�~�g���b;#K8��e"�S`����wz�DT�~q1`�����$�Ϥ�p/��\Y�Ž0�k��%��/��ebBQ��p�8�!(�>�	�X;&ۙ��>� z��1��A�!.��+�>%8 V�{x���Ϝ,�+�Y�r�6f�e�i�&F�J��b�^Z��P$��G�U�p�/2e�z!O�I��j;Z�%��ͱ�"��U^~3����}G�'v��>T�K�s��@)�<��U�+F�j��n���()1����z���<����]\�zq�9�|��SX@�;�����"0�f�J$(�jC�[x5���*�y�={(l�۸���������'�2Q�[�xG��5T��e�q�U��k�^�j���b.$0�e(�T�S���`Ϟ��ˮ[����l���޺F`y*;�A�#)�,!Iֺ����:����c�x�$&�,�U\8���|}P ��ABl����I:B�[*�ħ,a���!n2��4='i��4k~d�!\1d�NQ�+�LLRxQ�f�3ȭ��v!��mSo�ާ-� �.ne��MO���خ-�;��˥�j�ù�η�fм���L��9��/L^/�Z3��1{J��1D�D� � �����3���+1yA���������a2�73lgw@��l����F��ۊ�Kܙ�� �A�I,i���*Z��;4���p�Ձ���Ӛ�'�&�e�hy��i�������~���Dn\�M3�����]BK���H���b����Eeӌ?���Lц@�#�92��: ��XK8*��f�\m��Nz���0��2:��K�%e�nL�x��.�Za�J�"xbm�w2��4[��3R��CʔoS<�q�:�z��^�~Y/�Rny�~��n�t��@
�[�ui,� o=�z{�̞UA'+,F3z��ӾgŇ�����ΫƊ��$IP�c*����~$_���AV�W)��N�H�w��i	u	�� �`^ı�ϋ��r�(�Y8���P-_1�-��?8c��N�R%K��
do�n:*��ܝr��6p��� �Υ�0c�L�������T�b
{@�Z������'�"G�"��R:lm��1��_$�z���-����v� ����En��{A_,RG��R�h��+cq�!�q?s�i����g[�:&�#���y۩�@EXZ-��;�W
�QY�o���?9���-���/�Pؾ��RA�9 7X�Ⱥ�-&u���U�1O��a�O1�&;��r���\ޏ�U���U�����lDDQ�3Ƕ�l�}t �=���#/ Vt0˚KR���4�k��]���S&����,��E��_:+�t�+f{)ZZ@���5�W�e�y�ʃ`��G�9]I���Ϋa�c�:�eO�?}z�F��	�x��.�ǝ�S^c�G�{��J4<�u��`ux 4�����^"�"59A��˸|~�{ %���ռ��]c�L���f�I!�T��
�C0�dN;���I����.�x��e�?^oyRbRn0kk*6|�=T���*^vKQy�N&BiY+��?9�*��^���]V�m(菏ߞ�'bX��z�^;��zU�O��R'c����j���z��.к�7���P_,*ͺ�=�}��5�}���D�����D��Ӛ�����I���[
�ݴ�Q���O��/){�;y�(]l�sS�)9\t�[C�[� ����^����V��ԃ�O�}���l�0�v��\��������x�|��H�ja�6��væ�^*�נ�=�C�Ъ̩E%E�u)E*_�}��7�}l�')�ܓ�n7?�Rnq�aP�5�q�{�f��7܋�9 Ie�1\�&ʒD�4�;t\!e�a�QʝR~�צ%�b9Vؕ/N����/e�i �[[݄��Tu7�$��<�S%-��OD�}#F�����GX���$g�B�a�n	��� ����2;�Ĕ��+����*N ;���(�C�;��r1�V��k0T����z��hi�/��z�F���QP$��yw0��3ۋ:4�J�:�h�Y�JUfG�
?�r;KdƲI��������
��]��s�I���V����_�L��|�i�o��8��+;['��g���ZtD��4�ymyx����(\n	���z�o��8v����u����_x}�.�y����ivMgߜL�I�\���v��rh�K�J�S>�aLYo#ɮ]Q���qv~�X��lM���7��	z��kx"�8��������)F���h��n[������e��rIv`|a��H�pɶ^w���$���EFS�7<D�}�Y�s׵_����I�)m�kDm.TYE�!��#)��σ R/ ��	Ȧ�����O��$��
]"�UV�f�6Tp�Vu�3Ċ<{�
�����C@)J&�V3^Nt�Z0&Z�R�~["S)���'m6��eI�U���DŅ��ZA��6�HC�%�ӓ���o��RԴ��߲Ą�%�z���ftăW�`j�!e�T���\� �pL#w}�M�.2�ȩF�0��h�cиQ��#w�5���[L��$�0+�,&c�X��l�`}O�fE�Z��H��`�e��=�ݻY<\�W_��R):�b�M	�k������v�m� ÜM�C�o��9��{+�=&Q��?Rlf��	8	���l3~�_Y�"�����=țt�I,��x���8��R�D�M�h� ��s�BO7/�~  ����j��\\+�gN��?|��n=�/���˺�7*�z;Qk�uf���gm-�^L���i��M�X�k��U��#
�։/ �a��1ց��	�q��s�VH�X���b��V�Il3CEޯf��Y	<D;��,��+����ZS
��{E�6�!3,�/w���y���@ח��{3�<�R}f�p �捀1���gV�A����
� �����[�e� (�}�ʖq��Lq_��>VB"A��D�K%k �9c������|c�\����ag2�������`�$H֣S���8�l��gT:j0�P��R6*�/YRS�!!�� C={�}��6$7�S�Sي��+����iJ��X��𣰱�j�3�%�}��yKd�،㼠�ǎ�-�yK4�b����F�ג���oV !"�����pt<ù�^�)5�٬y!�p��Z��<�B����ґ��KJV��s;t����D�%�'<j�渋Y�/(�N����\.�Z�پ��~�آd��X�IV�X��g/)�6(���
KA7P�gs���]j0��(]�t9�UoJ���R+��6'���t�@��	)F>zdb�v,
��ѯJAY�,�5RT�ϼN�;����QzPV�h��b�5*H�G��K]#��ˇ����Rv�Ӏ�����ս��*�GzeN;%�G��e��橵��������Ĵ�G��)�F <2���%������"WFo����?Z1�1����_�J�=y�'��p��l�f@�nL~ ۺ~
��&G{տ��/��xj����!N�������ۻ��/@yE�5�hbht�E�|K��L�������PYѰ�=�J�I�@o�cL`�r8�#ǑYC�3�8��1\QE��w=���K˕^�z�ɜ��j���q(���sڊi��UOU#�"R&�q��!��� w�l�vlMc�m�	�+.-��_)2�W�4�f�`0�M�3P�UªXÆ<���){t}�R���<�W=b2Ĺ��5����u�e�	ځ�T�L�`��0����Ϝ����� �����!3s;�&Er�Pu�O��Q��Uv���E�_��#ş7Ū�+n�}c�5���_.ieJ���0�v���))�Y�K��S�m����S�i�(�Y��z�[�'�]��#����J�X>	��V�E]��	������+�Ǝ/6V�l� ��);b�{?�g�O^�'��[���.�R����X�L��� ���O�ؑ@�R<%`��M�b�@�+���@�_����BY�7C�	���q�6'�~q�[A�8a�S�W��n��}�{���;}cr�#�Ht�W�]ek��ʘ��{~>H1�T��A�T��f;T��V������^h������r�,7��)��=���a��:�k0֘��@[������^Z�@���j�'�}��d���z&�?G��}]���g���j������g̥�1w*%��%*,I���ݼ;�~�F�a�p�����������ܶ�KP��4�䔙�`n�
�*cV��T_|���ʪ��<���p��3t� l���E���\�V
B2fdXHu��?6>��ƍ���9]��Zg�ː�Of�}������D-����'	���J�~KE@=���mr��i��QhY���gSh��M��o}R�N�隮@�V۽�n�M�:\Z�}U�+іة1��дϯ����Y ',���_��T�bC[PAI$���޶��1�i� qҸ����n���®]�����4+�cX�����`���#o�^qX<|=�8ؼ��mO�\��B,<N4DH&�^�ǓIB���3+Nk�e��!cM��b&q7��_�ҙ��Pm�ǙM�� ���_~m�42��MP}7 ���2��a�i�s;�) V��c�t���S�5�<^ȋ~;���v�F�p5JhY�굚��c��ȓ�fjȪ��������� �e=u�ׇ9�~��3���i�o��̈���>Z����$���N9�"�	%��6b��\]I�o��?���p쵨��Ҙ��x��*���b�W�%�k֍����s��O�̱�T?���cPB�5X����ZAX��!��hm֑�r�QA��z���w�U� w��������ջi"p�e�UmWM *k��P$�]6DA��W�h�Ћ��U#o'3RW	`<�9�����%��IQ*��;�m�����A�5�Y����X
��Ot�Ot�pI~ib�UE���'�/o�u���=�Z�~��Vb:K���3	�7܂?�tyR��.��@�.�	 ��#�7A5;=
Ac��7�\�����[������E�����W_�.-[�/�9O�L1�Ͳ�H��R9�PէQE�2�I�[M�a+q�n��F~�Q�fZ+ޗ=g���@4��3��
(�`o�-��u�f�u���~����$���~�.�������Y��p�a߂tN̲<\�_�ѫ��B��P��*�i�3��%D�BzQ���W!W1��C�^��a>�Pڦ�',^X０��2�A��K����n<𐀮s��b$5�?�=����'��5?�ߴ���Ŏ2�&72�ة��ۓ�j�bD�Z�g�0��X���T�y�o2'կ�-���A
����So4 �e��*VV}�+x�9hQ^���C^��"�d1��R��lEz��%�;�Y�̯�(��Վ_Wq��r>~p  ޣJ���_'f�8�ӦC�a�2����`��&�"�rf�����'(`��蘭��Z��J)���U�M�
?]_ ie����)�������W7=v�TB��57����O��� &�Ꭿ���[�"�o��A;9��矅����&���o�S� %���\��Y@�|'B<�����D� ~�y�iSc�Rb�)`">j݇eUB=V�q������to+nr�g_A0ώ7�Z�$ �����G�3��fOt}����!����-�d�-�.���`�,o(�g�3\�Z8�
!�V���A'\0��-�&!���.Њ2�1�퓮o]KY`��寿��3�fJN w��4��0�8/T���P����;N�x�m��pGCH�{o�r8�̬���H!a���x���M�?_뎅�.�Ʋd�^B��~�#U�>.��rVp1������d�����
$����s!]�;L����Q&����E�k����@ ᎾÍQ
~�ʓ*��Cy>6ձ����	F����UΊK����1e�\���F�Ls���������la d ��v�,��.��f�6��f��ﳀ��O��7Q�@[@7Y_>�^���f�(�.�o�XQ-�XE:sz<o~%�D���Z�/�ի��b�gD�~�M�;����?�݉ߣ���2��g���2��0\�Y�7w�θ����z��ߌ7p���6����V- !1�������p�FOpv.@�"�.Y�o�&V=�"�~��i��
W��F��~0FTv񟂜 V��m�Eb/�����,�&k�4�Aҟ2�%S �?m'�o� 	!�	Ѱzq��wby�u�M]�p=e�E1��n�[��zeט'�X��f��h���ۋ��rz�㷱
u&��ߛ@<)�)_\�,߈31c���ˀ�jϨ��2*9�D��BQ�2/8݈�-��L&�H�Y
qQ��P3�դ(3���n��gL���J64jz����2�Kn�'��u�o� �%�߄m�+�ϫ�pn7c�ɵ�!�61{�IT�e�e�s��fe�v��#�P̈́N�:�s��Z?`,��=���~m��&p��y�l4T�����I�*�8�8(��R޵��8Sn?v��ּD����l�.�I�4A]WP�Ǉ�D�Ȫ*�斏�X�K��0�?�/��q
V�j0����j����Z"����^t*�8����zY?�z���+p4"<�S�����>)A�N�F�͡�"k��<��%�.�CST:o:);�r:p׀*�S,�^�g�%��@0	�#
M��ӭ}R�ˌ���u���k#�D��+��%^��|�O�/���SZ&�d[�U�C$��
Pm�Ҷ�Gz�}��(�ym0��Ċ��ɥ=u+���LwrRb��|[B����C�|K��4�(����D�}d:"�e���z�[V�P~-����[�eI��ۓ�X�$�����?h�����l��^`�VN� ~r�&7x���{c�V�4 ��ei�ؾ�G0[9�PW��'�bp5�(B�N�GY�-�