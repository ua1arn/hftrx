��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga�u+mq���ĤF�s��	�o 褲�[�P+�2�4cA^�������>�F�,0{6{G��X��Z��U��5 N{��#�?�$�}�eG��'�@������ff�� =5�P�TY01�D�5��# ���|�Z�T�2�ʻ�5�3�^՜RHK�P�Pp�餑�)�&4hQ���1���o��K}v��ܚ�[Y�Wv+j� =������h�%>�<)�	"V�3fe�5n�m�	(�t1�t!Sd4�����/��ЗN@_g�ν�mc�0��Z{Ж�-�� Q�BT9Q��]1ڱ�*A�v���[���0Im���=A�lY}��Շ�12��#t��m�8�N�|�9���T��l��Pմ��׺p�D�;\s�8[|_��	a�A>rW�#ȡ�{�������x��V_Q��#u+!�8Fm`����O��:'tS�G>bKJ�O_�k��R��#�Ơ�>[ló��y����54rf�� ؙ��U����Rm�U��ic��R6Hb�xZ]�ǔJ�Q��9�Y�J��i�bl�[�G4Zo�"�d�=�j#�����Q�n<�4
��Eo���Le(����	d�J��h�Q�I��2����O^���<h|��ߟ�i�5�ǀ�� )��ͲVίƓ��<��C{�A�z4���^�j��~JV� &�#�"L�ʯ��ʜ��p�>����;� p{ssd:y���ZjWk��]�}��ָr��P!~O(<p���K��j:��2�$F!�Ϸ���	���d�����_9?�=�M��5�>��e�o�`vп�����8����	/�� �2�k�	x_/��惝�"I�7��w���)7m��nZ�֗s���N0�YH��H{0D�G�4���.c��ղ��{��3J	lO��w1�ȓ9�3�7���VzV�Fx��kw�8�,&��J5V������
t����	�(�*�-��e����S5<!_�iK�s��La�ݸ�'߁��&�]��bx@����=�����B_���-��^{�%S֔�F�3ND�T��.Ա.Q�&SZ�N2�As��M��;��X�ϋ�v�h~�;}g�����[%�<�lƋ y�"���˳p]E�kTŊ5�:I࿥©�_���}[��Ȣ�"��.��;	RFƱUz+�yrd�2�:�-#��3~���r�΀yW�5Wa�ɛc�YX��}{Y���8�����>� �磰q��T�c�^ѭ��(�)q*B��	4~;Xήpc@98ؕ��Kr��o,� �ov��@炙6H/�d]�L8X[�9��h��p����4�R!k
���|����i����"tʅ�8$�*�c�=�H�o�������5�>e/�,�i�I�6!`��
:7%�F�Zw9�/a�*��K��$���G��1�(�/�.�ʨX���`1�\��L�+�@�N�*r)�j��D�xL�+}���/�D�%�6:�
al�E���)g/Q�܂�.��u������]�ז-s�GԿզ��us�$y�of����x*D}]1���Î�H�G���5�����r|�I7��c�w�X��?O���z��p1���hL��tT]�?{���(�7������傧������P �'��	v�)���V,�:�bה�`�H2J-.Q8:��'��(�L\�7ė��4��c/e�yw���0I���21�;���M��d�&,1�0�y8��}���4��t�QKa:�|y�@���[<S~C9�Y�����]�
b{J��0m�g�(Z������l3�4oL�kE6ŹS9%k���|�B㾣������A����0c6�\��R�l���C\S%s��O�t����y&�q)+9H�5�������Ceg��P��, �q��w��Q ����1�R urUM�#�A[&�%g��u�g��T�A;0Yf� �U�+������x���jVK@�������_��B�������/��K����wa����`<l��_���$����ЋMmp���E4m��ǲ�����<R(�<����϶����d�Vu�ԍ��Q�����\Ç�s�����<�+rC�%,�/g��Zԗ�D�iB�xY/�t�.��0d��t�s<�6 �a�3�"��$;�	�­k��T�d��{L\�F
�>S����S����H�M/tu�_��V_6m��hk[u|g��.��/r�n El?�1{לz.|fC���&���d�"�%g�%)&�[y�+��Q qz�?|:�>r���$�E]~�O���V�*�W�ҽ���K�.�4r&T�ӂ��W�D���s�D��CR��C�S@�R����uLt�B�f5O��!e6�mk_ZS����| �����Ek������"�5m�6ݓCfa4�p�#.��K7�7M��-��D~1:DT<��|"�!C�Ă��}����g�ʁ88@�0��� �\E�QI#--��d*�B�+n�a>��<eD��s���l��^�`?4�@���SM�PW�o� ���iuZ�B��"Un4�ԭ�[��Fi?��9�6�=��G^.�?��(7�?I�Y;O��)'T���2����B?W�]�p�����.;Kܻ����s)ݝ=��n���hqC[�4�8f�M!����zf�_���û�/�W]������Pf���J���{X\9B#k�u?˽߬��<(����"�ڝ�v�>���ρu�� ����+r���<�β)�/��L�H�VU5���?1��4N�z7*I�hG~&R�9鴭�<|�ָ(����E_���}�rޚy_��ؐ�i~󈍮Jb�"�|"4t����m��	�����7Z�R����V��Җ�v�f�K-�jl�1*0������8�0`���g&��D!��VA�g��󶦇�F��B�љpy��/�Ժ �.Aq�"*��W�a� ������50N��J�IȻ)��8*�B�R�H��B>�"��yk���	a���#O�0
<jɊ��׍�ܥ��&%b��&Rs{	d��7�A̮����UZ0��
�l&6�I���Z�Wʬ�!��k(z:9pWZ�� t�P䰥�87r�B:�¡Lކ���xO�BgH��GmUX����7�i�h�Ŗ�@'���Z(�r���A���b�Ye+���u*P_�±�����l�@l�s�X����'�l��l��\��*('@)�
���&�yB`"�E�ʅ�"?=�n��&���h��A��F~�.�!G�Y�߭�yٶx�l䞓�5�l�
�Ή��qpr���)}�_'�����p������/��)�wH�H��[��Z��ĈJʥ�O��
{
�KLt�m�p6�!l��H@�ŏ�>U��D&��L�#_�;�M��H��ұ��0P�,��K�1̈�BQ�����l!�+�ҽ�T��J7�N�
�լ��td�$�+��bw0}�\�Z/�hȊ3��&WH�6+t���a�䶘p�`��>%l%7�޴P=��	�=�>_�'[��U��,!Q�b�c��rn#4(��>=�J���ƞGx����*���nh�7n��U��x��U�%_�~�V���u�9�[���E�+n�t�x`�����p$��d�y-�OB��]Z�!8bg�1+fXFW����:�cӳU�{�!L��u=������Ӻ��yY	4k9��Պ�JV�q����5��b`�yo��}֮�y��`��u�&H˞k�לG�1�feEMuN[���g���ݾA�i7��g�y�
s��m��:��m�b����}P��U�n.�U��D0�7;Eh,iTr�t�<W�G�.�Ԓ跰s#H5V���� M����ڔ�m�_�2�@~]V��8�׆�S��>Rx# ��ﴶ��x#��q�#>�� �h�mG�M2��X� <�Z�)=i���ȿ5�$G ((u�)�1d�]v$V<�����綟i7IxpVq%a}BzZ�[�q�$o?��.�@3���zN1���4�V�7�Ίڦ$/"��@�d�[���k4�)X ֦�~�Q�����ar�n��8��m �O�6�+1��d�n#�D+@��M���О�(-p�������
���l{|D��aF �r�so�gG�	SD<��xh���t�� .Y����ƣ�#�:f����6�Ǜ%.���m���gK/�
A&i���U�x���%��t���69�Dh�=��;�s��}G���uJm0�=P��c�1��d�,�&Of��P�J剴Z�܅.�Q��6�|F�3��!{�+��t��Ż��z3%n? ���xi0�ĩ!{��pH�P�:�:�^E=��g{Q��9�ÚB��Cz���O�v�S\jq�߅��	{&C4���'��Xe6�ܟм���
�Xb��KM����NX|a��JH�	˿t.
po�-���c�ۡE���w���x�eu�l	�~�[E�0K,�������p���h�мRw�OO��X[�i,�ɨϲa��*�_8�� �XhɊc{$�˵��h��D"dA<H2&�#�b��#�9d)�}�݆����&w�UY�~��6��Tr�5ؤY�@��R��m��@A�o�zH����pP��,V�8���5��������� pf%����AVrT��RY�3��C����>s�[��3�rj��).�2#��x�eR�ĉ	,Cw3�����ȯP����!`Y��~j�9A�=�߉QN��#�W�����+��`��i4�@��@���0�)�ݓф��=~�C��S�ѷ# P.����E���(�"�.�R����\Xm��~,o8�,��=W�Nt�Ƭ�"�@M(K��O{��vHG_���%�����3`o4T0dgвD<n�H�]���e���,�k�Y�(��m��r	��{�t�x���K�q2})�U������W\��9s6�����18���'[B퐲��J�F0���1-\�]	�6���=Ie;��^X׍ ��s.�!=�����ñ<�T����(ugd��q�	`e.�N��i�2l�p"39����d��1�w���IO���)�1�	�M�"���;�v�xo�Ƴ#��Dl�A�d���������j*�<]ð���Pl�[0�sb5R]�{>�}���=wwO�&����J⣟��C�Jn�J�ϡ���������u;@���w�	��C��[�s�~�GGi2��k����ʚ��q@B)7�C����΍�}���]��'�1n�0��(3#�H�H8B�c�+���W<-3�Ht{�/�G�&7�wЌ0�%t	D��N�Q���tl���_M�=J�`gR�Ŗ�^�\&����>��l�����{��n��ڈ�%���̭U�rc�h'�d��bNz��QfhZ�J�!VX��.E,�3C7xg^ϚTS_{H@��7Y���__�����ŏ�ZpH�� o2$�h���|!��~�h�T�.���[v�q��^���~X���q��/>��w��g�D͎���<��'����;�����}������7����$R�U֡����3%
9�7黍�^�pTbm���r:p�e�Az&����1L9ӓ� !����M������6�t���=%���|ق�������	��> -�P�C�.5䔋e���-�{����uSɄi��:��~��dN�L&Y�qw�sM��(H�5@VXU����z�S��nܕ���A�f�}\=�|�`~4cmW��޻���U���d�`�is`�Y9����� ���۰��x0�w$�j����������9+p�ƠX�z]��uA�/�������3D?�M��IU�.��-��$V�W�Vk\OkN�H�t^>O��p'�߀	�y�I]�@��8�O��> �x� |�gcd��;?�{c�p�Ǖ���,a�Eh���[���,�ߒ���A��f���y��$����UEs"��S����=�Rv>a6׎�ҊI��W��h����(�b�U���+춺���Y���+�e��;�u�H��s.�f��!S�fxǨ����	��/��`t���`�P���^K�?@r�Kj�~G����39���4��[���26M�ya�N	���Jօ BVj$��	��~S>u��5�K.Ɋ�k%�]��Yg��S�������[�	��˭,Xnb�ܽ�Q:Y��O��J���Yv��1.d����/a7Clb�7�Hst ���w���rk�������Ie��Y)�D0�����*�J�����~�lr�胋v�E����+<����vd��֖4�g���V�1H�{U�[tf����Mkw��]���V7�X�����qT �Z��"��ks*�Y�E�@��k����3뇂	�v��\}8����l���x���9s�Ұʌ��� ���n�t�a�+�W��#+�ǢfY�(Rٵ?��i�f�O��8�b�$mT���@��L� ��:�U�p��㋿<m�DD7@c������Q�1|�.t����ʰ�W�o��r��Y�9�Й�2�ۑK�A��č{��͟D��M��i)���g������c;����7��!��,�)?ؒ5�����Kj��ƞ�&��E��!�#Fv��|�&�&�gV��V��Iuب�f��4d;���:mVA3��?�=�,[�S/�4�C��=e����8�mP�)�����H�'ENMN�4����fאN���y�u��;����������	KD"��C6��_�e����j(-�va�o���7�W���tX�W�; �����y����.��1�6������.��k��1͓_ t�+��ar��3�����q����.Kɇs�|F�⋝�E1a�.��
�m�L�X���)�$ϭմ�؈�8����p}#�g$Z_��S<�v[1@��� 3�x���M	ʙ���\��Յa<'oz
��[ᴟ�;z@�*�~�W��>;\����T�L�Lx���a�לS}��jiW̐���+���M��<\�j}�2;�x8͵i3j�-)N���J�P�8���Ψ�A�j��6�`5|)'	�&�qb�A�͖�E���A�3���i����ha�M�j	�Oz�K�)Xpsپ'S��*��S�j5pD��Qu�1{���߭�!a-�$�N��jl��uMR��� P���(R6�w6.�yz5�+��� |�1Y5�b<��=\zi�M����8�E�����H�3I��j�M
|��ǭ��jr��g��mRuv��H�7�+�I�v,b�;�GѬ�؋��gb���?ܻ	���"y���]lt�B����s"S��>��gK��@�'Wp�՘|��0�-R7+�|]�ڳD�����j{��r|�C�Mf6�V�G���IZ���,�����Sx$�Յ����N�_*H��L��%3��������zӴ���&�z��A�#�k�a�W����ZA8w[`�Z8
{�P�k�Mճ���
5"��K6�o�:��Kv$�O"��v�J>���{T'T
���f�oh)k(|��g����ĵ�n�#	ى�[�ʭH% �0�4�S�i ��?�'���䞶f�����60����D�$�נ\����{M��`�F��O�2}�ZI�i���ݘ)q�krj���Wz0k\W��4��OS��Q�'�Л�Oټ���a�K$Pa	��ɺ<�]'�;��?�ʜ�ǰ��%S��%��l��R`��fi7��-��S%��,�zd=˲�~��ޠ�ʡ�LL��
��dz�0O�*]5�l �?�6@���+;���+!���)�Z���8�Zu���;W������䵕=m)ircn^��2��*B���6#$�v��lDd�\�ڶ8$ݨ���D��;�/-ת�]{r�\�dr�t���}�Ȝ�ٜiU�,h�:l�1�6}�l�'ₕH��@�"E���
��o��RB5���qC�	Bx�DK�{H�\�h\���"��zT��b��r:Ԡ$�#���V�_@��o�����J��ȟUx�J"AUAb	9 &e$��ym �����)��U�Z[��̴�1�'�
������P�|.���,B|��8�4�*�Z�u���m�����i�����5,����"��&	ΰ\Y@u��>��jb j����x���Pr�O�"3;��u�9!����2KV}��/��H�v�_@Bu�k��?o�[�7�"����A�0Q\�p)K������ZV6���й��܄̋]>Q�q�Ɣ�hH��;7��4�XG�$K�[���%���(��Nf���
be�X�~sa�I���kf�:텇���b�8^����pؗ3:����|��7\���������Ju�8l��1>�P��Ů�GxM�Y�r[��9|4o��Q����+�=��7�h�WϷ���&�4���,��I�|��	�V�Q�X��.�����:8�EI��t,�V
��
��C��7�ѕ}Ǒ��X&j�`Ԑ�7Z���E*�8U�0�xw+��3��{�!�7������䛢xQ�Ksf��P����u2�M4�����W^x��DU,ܒ��Y�i\�(Fܫi��1z<���a�Q� ��5[C[��/�OܒͩFO8{��Pc&�� ���^�]�s���Q�����޴�MR�i/]H�-A�!%�7yD!=�g�=�u��7\B[�F����U�Q^����LY��Ō�	6�T�}j�{ `)/���Pp�[�:K��Q�����2�p<{ذ���U�vU9��av�y }g#����pش���t]K��Q>�eVI#6 S!��a�k�f�Ï1黳$"�>37��V�(�;��j6>)y���Q���eǴ�欤y@Ƕ�ǧN&���Z{�M��M#�T����#|�i��!����2��dO��$�d��w&0����J�b�/k�X�D'R����o$�pM�l���&M��������TM�������yF��4�sֶ61I�'��B�L��Arfkv����l�}rat�8��o�6G�Hs=�;��N��o�q(�vࡱ�(���;4��Fp?Ζ�i����x�3@z�	+/�ԶWz8�y	Ֆ�
�^�� �>�^W�b���tئ.����EV�5O>
�]�/	�h���]J�G3���WA�ꨳ����M`��,�ĺ&�^������:Y�O��z�, s�=���4���ҩ�[$r�~��+�^�5r��U5�f�Z֟o0N��M�<ogFQC�q�;�
)X��6E޸>��w&�0�2�I^��:M���'�Q��ߚ���R:U�{t�}5m(Jy}u?��8���` g��oVp��!�}�����7;��b�K{Y��p�E=Y��ّSF���U���D��Dq�g��	�����F�#��ix}��Y��0��:�.N�G�UɅh�2ET�[ ��n�3S7�g��AQ֑�������e� :�����Թ���і�J�Óu��Z>_��WP�߱�e5�2���A�c�U(����u��{Cr�s�����Cs��|�9��)��%��-,�!���}2-��x���$ ��4U Fo�?/��Ԇ���SV:@�7�'wީ��j檎W��VԌf<��=���^��SVv�Z��/�#�c�vciwLN�q��om����<z:��C\�1} ����Y�6n-��k��t�W�Z��������e哮!ZJM��{@�֍5Q,�ن�ct�]�i�Q�?�cc��vV!:s)�^�+��}Ub�����ls9���n�֥i�d��a^��;����嬹4�z�3��퉕�(�F�'� �� �@������Ռp�^n�eK���V���X�.]R�h#P�1<hx�|��团"���6���^Ӎ@��!ޯ�a4!(>���M��-`P�H���&�������p�����^����N�V�D�P�x���%:Q��	*o.'���1��L�vB us<�հ�x1�Ub����/^���ɶ��FKF��"�/��ڍDa�B����<�S,���O�U,��%�"�J�M;M
A���r<�N�[�����q�������|BF?N���2�0���H<?���.������v슃pE��ڟ����dX�	��PG�5_Ғt ƕ�#�s1CIu,�f�f�E,#I�|�"�������k��0�dr��.�J��
��y�q����?���92�5��L�,�7�I{Ҽ�����H[��|�A�)���h�,�nު�6&�{�y�2�}�-1S5Ǻ=Z��[����k����S�f.�=�Li� �ާ�����qT�r1_��d�������q������ּ�K��!xM71�&(�=G��%8bn@I^�6!��̮k�-�3w��L�R0U�׌�1���f:�d�	�V[�w~d� 0�'>ϵ������ac��������/�mZP-K���lY�`B��zpB�pސX-͚�~��ӎs�;���ր��p����+H��ư���w��s�	8��E�)�����i]����*���l�Y�EF�M}׭x�{�
\�/���$�t0VΆ:ǫ�N�h)���}xޢ�F/}T�9F�.�+0i�c�����s�d�j���F�#WW���$z�e�iT����߂VCˎ»x��a�Z���D�^��ή7��'�_�P��_�W=�~7zX$�׌[^��W\|�`�6���9�Bӯ`>_�m�t(�����Ov(�1�st��<�����2��X�=�ੈYs���J���$ЮZ�f��ʈ����\D�#�����aK1��Y8������w��qU_��|���4��U�m�J�+��3u�/�ĮMz�������w�-K,�c�k�BM)7�x#A��#�OG�������&
�¾_>�D�A6{�����x�X��<�F`��oo6[�u{��W���A��S@lg�׹f2$Y�B)�|���P_��5��T/�udk���m�Hd�5�k��s�!APq�M����9r����e� ���ĥ�|�!@<�'\�i��!�|�,��\��@A���-"P<J[���M	|���WldkTCf:S�&�K���o� D~���T땲�aQ�����)Nr����m�	^狉R�,�x�F��;s�VUxcU׳c��>{q��_?e��hH�@��r�5(�;ٗ��t��X�A���˖[�c�����7�����)c�E5�����h����RF�+��s��h�Q����;EzE�Y�o嫈H��ڽO�Y�zOY����X��#nM3�>�^B���5^��s�8����(���6ވݤ�Z�s�h
!��-�vP�ʳ�` ��*��!e�\J"C���z�'����.4�j���4R2+�|67�%��26�U��~@h���^oM��n�
�2a�Bʥ�]��Pު{�J�E  ��y�Czp�� ��"�Ƿ��jL��X�*�!?��@>N�m�DҚ:�,�4Z�S���.M�{kI�Iy$�ֆ�cqFF�=�lܖ������$T�>��5U;���|�M��$�K]\��f�_������8n�=q�٢�Í�5
Q����4�1���sfB6h�zb��|�
b������KF�X�DfiF�g�����o���qI�A2�&MOE�x����8b�=���XPGUk^&1��]3rݖ`�h��� �_	�PeY��M+U-�������[8�j���j�31��|U��O��X��_1��t��
ve�?^$�*�(?��ke�������Ld����o}��Ǫ<4���<w�'���,Mڊ����>�i��(�@��=�R�QȈ��J���߹a{H�S��%,5��Sŀ����W��g��J�pA{0<�_�i�(��T6=�6�S�6��:}'�:����S�C2�'b̦}��X��<tzI�������ͦ�x�m�<��λ�xܰ�-��*J�}멹�ֹ�>�2��0wzZ<��j��L�MYY��f-��f#a�˅�^H�݄�e�:(��/�{���Y�E$?+^�ͩ:���hs )��;��?��tĺ�~�����^��\?a�^KѶ�g�As��'D�.��6�a	����f���T^�밇��!�>6y�or�S)<�˖eβ��N�n�؁p�n3P۩�,Doǖ�wx��=�i�U�Z��x�C4���u���rk3zY��7m���#cK���ϱ ���ܖ�=gN����K|G��J`=��`D��)�8BxG�Â�Є5n4`B��B��q���]r�6�յ��΀Z7�S3�qծھ��cW�s�ZGI0�N롯��W&`�o ���wZ��gݑ|봂E��O\��7/>���"`$q@}�	���,uj� }����F )��=��a(�Ў�vO-
��7Q�qiph~�&����=��dt�ӕfk�5�� ��4�@5�;L�o[M:����nh��v-�t�%Ԛ���f���g��$.��S��Lwe�r꘨���Tys�b�l�7�G,U�y�Z �bv�T�]}T�&L���E���9V��ռ]��e۝��gh � �ȷA�,�>A�[���$T]�/~+�j^oѕ���ˋn�S=Y;�h��-�D���Z��������	�[�a�&����g#�����O�	�yL�ע�:-~�M�۵�y��XI|<�୸u��	�� 5c�ҵ�?L� g����P��h��4d�t�r\F�h��S���lo�1�j�90�����>AJ\D|8%�����\ɳ,.�x!i�w�'�x�8XO�q{�S��N���7�H>8�:B�痬5���F�'о>KL[�t��V"�>c������w��2�IGu#i9�(G6�[����D�*���;� G&o�T�.�LOb^��Mt�l:�eQ�f�#���Z����s"\O��?�#�&��Њ=f�[�����U����Ѵp5'���GR����n$������*�U��/;��6pW����c�|"҈�14�+���Q���$��P*�װ��Ͷ�l����d�ΥMdUH�� _�����Ӥ[�F�%%�M���U�(.�^���WW�h�~����-< �w��l��}���(�mNa&�b�7��،eU#ƞ�:U�2�FN[�ђA�*�J��X�/T��o. �� �Ć�O���e�������] R\Ĭ���xE�y&�tb��y��}�ou��r�]%�ʃ���8�,�6E6�g��)0�mٜJ�$ʹ�f�	�N��Cl��>�_��+jI\=��"��(K,�fwۙ��d��^yJddpF`�SkMw�C}�8�?��-!�|kw�L��3�,�E��k�{����=�}��`�jd��A|�8IF��|��z5���z�U���ȻlU�������~m`nY:�����rY��cƴ���_�l��rĔ���|�K�a+�7��g������ج���g#4բ�[�-����(�o�3%���m�=���2Y-��n�?�X�5��&�j��T<7���Bk�~&p�L�a׹,<��2��� ρc��3OGRQ	����C8��z�ł�j�O����R�����ϰY�R�n��}�Q@��X� #�NNB�zvݕg�E�O���1/��@ ^����m�]�Z�������7�[_|t\<�tl��j.o���݇��Փ�������U��@���k"�>���'�Bm������D8��r����D�Mؙf���}�o/�<����&�	SQ��H��V�����{�{�&]�mP	,�>�����1�*Q��b��X��e4��2��}�t����,�i��b��e%�X��E©��՞���8k�i3�1!d��6��h�P�ۮ�Bp!�5F����r��|�k��R�¦?[7�VF�G@��'}��D:��y�i_�����q �(S�!�E��:�ֲ����'@�F����$R"ЊGB �lu<�>��{n	�vb�ڶ��]�W���K��ҨT��Rb9�|	k�����|�d+^^+B蒰s�#��񞋺��ݘ_��G�Ռ���qt6be�y ?�������Z����@ȅ3��d�� ���&�aW���t��LN(�<���[�������7�M�֗IS�c����\;����P�K� =$0��BNO[vOս����ǅ"�ۜ��o~�d�RX�!�%�"C1L���|X%�B�� ]o=�3=n�?��'��7�o/��9]6.c.)?u
ӡ]��Nd�|@g .Wm�2掖��S)�̎�egL�K)�>F1��K5̵��{�Nע�vW��(�	�i�`�$�n�� �äSB~.�0d��59�9�n�-���A_��G��"���!2:���WjX�
�X(�s����{���
����L��&���1�l��;����M��!*/�^7��Sۼ�m�0��u� �r0�2̭~���|f���>�-�����;?�W!�����|7m�$�I]���o��:~�3,��]����%Ѕ7�>V����X?0p,P3u%q�%'��)l&�
��UF'�D�`�5'<�ᵟD�K�I8
�`�9���b�p*�NYVc�(���I��m��䶊c~xQEMQ0!Z���&C�n��l�<��b��A��y��y@h\0�kI;i�w1��Z�H���^�����a	�9�#m/�s��"C���N�:�º�?�q��A�R+�W�!yW`uBPrK������co�ӌ/V_�׊s�[Nȅ:�@���h�C�"��M�k�O�X��j3�@����~�:���3����h-�����Mp�	��Ŷ�9�.�<�e��p����I��K<DN@N�k�3�C�@*J��k�=��gz���JYd���i��N��U��0Ce�`�F5�2{��V��8�݄˹��K4�-�ӎi��~����V��%�S�컆�����?Y��N�X��<��	C��ۉٟ(��̵Tk��%!�]���������G��˻^�Ym�66 r���埴�B������1�)��+xu@��P�P4�5O�t�o�W�s���$�_�WgDΒu+3��m����f�T����qn���@JFX��S��=`��Ԭ�Ƌez������+(��h畼���eM�K��#���T�;�5��(f��'���'�#��2��Ii�՜\��R]�6�����X�"Ez�?�����a Q.�N��~����L7�u%;�4f��\7�-���8PI�l�s&�eˤ��f������y��ZqT�] ��A�OEB�Bk)��W&I1;�z�`P���h��:���!Z�Od×�/�H샷�P��d'�G��ƌ_���%~��ᙁ��?�˿?�EB���@�}t>�Sq�_�-���]���(�ٍ��!=$�!��aU/�o��:&-�o܋����Uuu�u��*�Ko���x�X�c�������}�f�Rm׭\c{�'V����`VH�V�p�b�w2��@��%hA���i`6��`v��2��o��xg��O��2#�g ��n��N��|}$�"���-'��9�8ِ8�}a} C# -��T�ZyM���$ʸK���Rn��<�#���+c�%���i@���ƭ<+�	p�o�3SC�V����D�Q4��nI'#h;��R��u�΂t��\I�9; Q�E5�{*���]r�Y��u��o��/��
�����H��(�l1�^G Q&p��8��UlLc�
�tg�G����%�Am�]s�����8�W�:i⭿�n[� 9*�-/)����eT�('j��V�D�z���Db�H��HC1�����rN#F���.���U抒sB�E����N��$sI7���K��vp}kPK��Sf},ݬ�}C�s�	c �J��?��-��a�9��*+@+3�Q�r�!d�=R��n\5W�d�/<c���-|dun-,B�e*�x7�HpvՖ��pP���9�b
���3)w6uz��i�l�l�����_�u�!xA�����j�hv�ɮi�_ �A�O����?���Y�Uj='/ި0��`��0�|�u,p��!ѯվVkC7-�L�b���D.�lW�)L3��������=���8��g����{���-��"6ؒlX��,��Z˧���.-ŋ�I`��b�!�Xo���4�A�A�_�b� ����./f[�t��@z~�ǱU��Ԙ��DJu��A��~��<�pmش�i�/Q�@a6���!�h��à����9}�h>�ռy�k1��7{�k!��hY�gz�ϸ51����#%7����_Nl�41sn\:=�������_Z�+��:��P�ی����wm�*�e��o9I{��Ѻ���^���ek����HFi�cL=TF=i��"m��@�t#U�@�r�D�3l�L'*�*s��q:�gFU�%����e|��qZq�?><TdȮ����C�������&WTo�L���p�)�82l{���x~�����o�7u+��6S#ke3I=K*�6J ?O,r��`�~\�M�f����)�e���w�ZQ��I�2o��.����q_���.��=�̌S�7�o�����V��dN�H<j�jŊH������\���C����9�u4>2�����}����=�4�JCa�ouD�H.�k{�x�Th�e���Pz�ՎŚ^��k��b��B�DF	�b��3&��u���F�J�!��Ob��:�\]���51���I��\������Pb�2��^��v���PLT�G�NL8>&_3����3tr�M(m���R�@P�p<�T������ǵ*�lL<-U���G#�����j�V�O��KBl��
k�7�f�� ��>:>���Q��f�a&�Dw�P�T�lp\�}�ed���Ç��_:0K��y�@���6E/�4�k�-6q4\4h�,�B�;?&_��U�)��5��W����^����m�0(b?|�.���T�y ��{��n��G�، I,��2ߌ�Xy��;�> q���p9`v7�@t��xQPB9'yks���APχ�q��L>䱲XU��M-�G�6�r��]
p�������e�&!R�"�?ȦUR��D~51:V8��M!�gf�)��
��8���������B�atM�\w�1���x��kTՐ��JAg�a;%p=���C�ک@���?��&5?��~���j'/� V�e\h%���忉�{��#8m)�_�U���O��j��Y\��z8��U������l)��`�_
�@����b݀� ��:D�[�|K.MP#UƏ� o�!�e�Ѡ�Xo�����^T��?s�;>��c�'/��s.���<��΋nS�����`�� G��A0��3���x"�N�09�M�Կ�×��ԏ�r��h��!�ETٵO�"�+�B��4�E�)�ە�G���t�?(T�T�y����Rq�-N��j/����ͧZ&��]}�K23}Bˊ��C` �!�O	��Dգ�kC���'w�)���Z��̮4������ʭ�u�X]De$�yӍ@J�Y��說�l�6D��׳7�Æ|B	v>�w�|�,h�6Mx���c�����i
pW�KK.�{��n�mw4���y����ܶ���S&��ᬌ;V)�u�`z����6B1��l��r7����y�-2XUa��zX��ga'1�v�8���}v��v��������y�[�b��k�,�+"��ui`r��bŌ�Eڍ󷘘�ps�b~ 2��x	�5ָ��e�j��a'�:��k�j��z�6&W���=5�E�\}����4�,ݏ��C�8�9;�r��eZ�+](��9Aum�d��e��7s��$�L�z�SzB0e�b��}��2�m;�;��a ���(�ȇ	D����-���k.�ckS-�T�=ߡ�[e��
%����	�_�<}�\�{`8m���;�;C���+���S��ߟ�#G��q�V^���$4��
A \�RJ<�54{�E����?ֿp�q��v����ll�{�dt�?lFK���{����J�`��dAk_���D8)�7��,���J�6�hW�7�Ѷ���g������Sӄ��O)R�OVq�I܎sL��<f˱�!��2bpʵJ>�@�j�j8�2�gU/S�nʣ�U'!sV�^y�SXR�&"c��)���^�!՝�︛ԩ,!��ۼu�X�S�P4Ɏ�P��͉A�&���\b���dXq�<}�8��P���RлI
��U>WRn�;/�s��uwS�0�����?��V`'��M���#uu�:���dY籒}ޮ�9��j�㻗�?�i���JQ�]_54� �F*l	��(���~�3�Y�+cz�isF�詪������XDh�-I�A�9O*��J	��|@D�8��L�Pn7QݔNmiw0�+�x#�$������ L�	Ȅ��۳�ø�����;���ɘu�Mn��E<��T��L�����S R\w.����e��kk�Ȕl65�i�<*`jU�N�cK�.}
E����Ԍ�-� ��
bXM;kzO�P�vh��k����Za��r���G5�G��S�HƐr��.W�&��WMڂs�E�
��ufϔ1��'���r����.:.~#�g�DU$19ݪ���g���Q���o��_0x�;��F�S�5��7��پ����+���G�	��d�V>ᾜ�,�� }W؂C�����/ ��FS^=:\��_\�/ �b<�%�c�{�^����4ͼ�`PbLY�َ�ę_]5��V�i�d�W쉃@��Ǥ��(S>54�&�>�x����4*��֦f]g��S+Eas"�B:�"̠`V�Xث�� �dn�m��,2����vW#�z��m�ZS���r�wӛ#��M�u�e]MJ�7Aq�p�/�#�ՎO."��wPQq�G�5 K(��ya�R�1h���J1K�Mp����s�`$�B-��Z�S@8�^փ-*��I��>�~D'�VW=�F2k]�J++hޖa>�|���q�XL��������A�!\[NA2�J�8�1+0ޖ�������K�O���ZD�q؋;(��8`؝&��
FIhK|V�c��p��k�]�[ԃ���IN{6����lѭ_TF��fFs��
I��s����&�)�����'��0=�Y�-B�S!!���~�n?Ό@4��zM��iUFxS/��'p��R����M�2`Q�2o6ޕ��QF7*4E�%���b��,"(��2�%|��Ez���j������Q�A�F�0 ��D%��R�iI&ׁi4%1�K��j	M�.{�#p�Dx���Q�A��韂4KnzDkߴ�-��̟w��c2��o&�����r&�c�Yt�u3OQXG[S��56�j��g�o&��9�9 �AM��kC�n�aX��V�l��t �ϘE��a.i�~�o�%�l4��e�Pc;��G�JҦ�R!a#Ț�s�g���n{Tq�ʐ�G�� -I`�L�8�+�o,wp���v�*3({?�o	��2����'F�j(�F{���"}�����B�Q��l��u�������òܽt�163��M��N�yMe�{̑�v��w��T{'����;�����F5C���0��)�L�#$�(���{�1:~�.�U�
�JTu
]�NQ u������J���Q�ɡ���첃LhB���q�l��BB��E�|�5���p��ZiV�Bt�%Ǒ��V.O�c/3����C �b���P>�}�S�/\�sһ��׳���03�9v[5&�v�{P���<�� �v철(��N�M����AL4��"�T�M�t��
%"�'�ײļ�j�P�g�h��;�ej�k5�����:PK?n�g��`x����"F�)�`�-��>-��d��@��g��CR�c������r�S�϶���˷�
��'	9ǫ���ʴQ9z��(Tc�A�-����T��.}��D<=���$�2~O�����g}d�A[�i�?E�I,/Mm`���-r͠WP�Bd������@*�����!Q_v����l!"����:(�L�+�@��Hy
G\�HA�7���ܸ�:s��Ct_vl}Y��=Q��(�7F���X��3�G�� r$S̓�o�r����(�0O���_m�F,�VeCT����!����Q�8M:�Xֳ1x�g���m^�����M? +}�#��������Y��BR�򝪍t��<��^7�uǢ.���p^�R�VfP¸��y��D��0�(�*\�V�/��[`9U%'kR����d$��E�enȈ,Ԯ��v_"��|���4��׿�`?�������Ֆ�*g/����v����hn}�R^��#L?V&�M�n�ĢY
��'bVoaB#F��H��T�*9F�i���s�T��g��S����]8W�7�a��v�V����y�!���ҳt) ��9񻥘�wÅ}kkQ��|ԍ����l>.��N3��;+aQ����ږ�7{��V?�� ��4�(�J��Nf�O�F���Ãk��}� f1R�����[����k	�! h���þ�Dﯺ�]�oS�	u�Ps�˓�&��ŉ���׶*>m/�>��J�m
��Ȯɋ�L� �!8 k&ؓQ��Ҷ^*�7��_�����0�8��U�[f��N�dE>1�.���,,<x#�k��$g)XnE��B�e�͐��b>��U�?�Y�Dr�ʟ���j�&J�q���$��1D֘
��7b\�/����n��`����K��������ZOM*޿���������cA4cP�����\Kj�4�e��g1��c�0���t$�!݋[��A���JOHCei��X�j����O֌��I�����rk"���D�=T��Z2c��]T�fl�Bk�(��}DS�e3�*���bQ�'��CZ�`�8�$o�*�ց�̅$��1�y�
L
�h��5F�.d�ě66�3rk�sJ8a?�0݆���%�.���AшN{��^����x��0|ʘ�$3���ddEE۫�TF:��lh8a/lH�5 �j̝���e��',��]J�����^��j�Ws��[�ֻ��m:Ӳ�����jJ!��ъsHr���!w��z5C�[FcV�!��xoo�PN��p�w�0Yet�QEO�#t��}��Eo��{a�{������MA;���歷Duwf�S�<0O.���\�g�J�ۧ*�2'	\W���%�9z"K���������=mTub�uE��R�Ә��_���k$Y�z�o����M}q��hEL�e�/Y��K�Z�9�b�G�#P�t2�S �����1'DF��^n�'B8M����іUg�\o��w2�P�n���˭�Y�����z��Q��6+A�2���T�Ό�r���]��s7z��4�?E��QD��㖻���>�P�� QK��>��JE`#�� �5U@og��$�il�f���Y�
��*��=g
L��h���{�g��"��X��܌�d������úu	Q*���!�!��&7��`�t☺[J��5������2��漘?��62V{/�{�S�is�Dr��L6y�ɣ郿4�{jbW�ۋ�u. }�5�p
0@-�7^�u�N��K>a���n�tO"�b�������?rh����;����}����'��d��c�w� �O�@�kz@`8s��7:�d���{�E�iA��M�����K����V�����%�1U�cn��!=���>�8�=�7�� '��5������vn�����n�ɚ��/丅���VK�f�^��'\<\�§�N�s|`(e ����Y�6Y��8�x�p��mNp }�f�ҳ�����Z�۔gƱ����ժ]�
?o1)� =�P?��]�8���6�%��Hާ6H+vtKr��g^�E�b�<(�4�*b/!ڰ�
��^��B��4/����H�Bl���������#�z�����<�ִ��s2���㗄G�V����c�S�p�E�hW:`�>E#@�������B��o�ƞ��l�i��3��)'����}j���	�X��V�ܡM��������o�����ү�C)��'�����C�Ñ©I8���4���K��p�4��🹗���=[��R��4���F���x;!çR�g�0%|��J�d/4���<W5�ӥ+��p�ɛ����Qo<;����Dޮ�.���+y��#�P�}�:���OWօ'ko��r�����<�&�d[��a0�7N}�J�6��I�����;��F[���$U�z9������f��* 2wϮ(�H���eS@��%9l'�Mل~v؝�V!�A��Գ�Wa�,�YL�fo JQ��hܷ>i��1�
wVG,0��V�N �	rg*(s�51qJ��%�h-�B�؞4�y�
����v֐�b}T�I
����8��/�(=7��.N!�['�IO�
�����2��b	��W�|������g2�3%Ai���l̀�?���N0���L�����9tz#�:� ��QY$:y�C�:�{��-����1-���J򍆕�a¯�`�D#(�]���K�����Jw�P������Ye�X����؃G�J,%���SW+莎c q�$�^�7BX;�~��8�-[�&U�P�9H��%oբÎ�B��j�y@�����O��@I�΅ۏ�s�L�X�܃�~;ΫI�"Kұ,����Xs�����SfKyTo�� �E1�Ju�ܔ�lcM��G3|
������� F����O
��W��F ���{"�n�`�+2<��H�W�h���$d�ȴ=���W(�.����`/2O���� ������4(���]��}�$�Xzgv	"�+��U�p-�گ�zV�:���"�<c-���m �(�B0u����S,�Q�B�2kҝ��ج�t�c'[����Jɦt�E��#� ��(��Z@�8B٥�y�b6���z�;��좏���k�h��j�2���g�D�
�Z:�ܥ�Ûp��!NbN��`���h�T>g�X�򯳹sZ&�_�����9Ü��&Y$(��I;$_x����-�q"�4u�>O��A߿�l���ed�{y�zi3�(�߉�UX�B�J�n.B��r��ѝw<��^=��W��	ٗ�6��]˼��sawE/֦����G�W[_��y>�%c�����s�ͮ��Ďj�;C���@�����-h����.��d�O�_��<t:�XƩ��B�SI�KjRW;$�.H�(ݩ�ړWq���<�(��1��W��:�}��V��<$i�e���~�Q3���0�̨�M�˲�2
�h�
n\cnnO"�w$!�K�}��9��'U���FD��@s!�!$>�[��zl����/�N��e�υ3��9��/��C�	&(�ɔuG�6_�����zO-HQ�DؽO?��f���"A*t6�65"�ݞ���|zn�%Q�~���X1���`dQ���Ao!W�+K��W���N��Tq�a������Ưqb�:������^�<�W��I&��aa�L��0ڨ	���YQc"��թ�xD��	�-�)Sm��i����z'����=Y��ɔʎ���_�x}��,�������N0�Ӎ�Q��ۺ ���	.@�B��vo�.�k��6��0/���.�ܟ��<��Zy�|b�[�=�n�A�sV{�B=aU���@ӈ�ڊ��|n�s�״�D�����.:���މ�E<(��.�<�D����8��zc~�Y�XD��^U�W��.+6���lP$
iŻ������ATr_����u����f�4���׭X~#�ο!���x���y1�S \�'�E4m�!�#����W�CbEv�z�`ka�W�Dl'HKS�#b���� ڮ3�~r��I;7���0���3������y��$���-b��,��21�1��d����%�J��7�+&)�#���U�/�@Y�������J�J���'h��[WJ6���c\�</��O�e��.<�q���.jF��;h#>S՗"�FV9���Z_�W��`�	��u#�������Lo�
��&<�#
�s�!�]9>0[�����e��n�d�s BZ��w�c0ݎ��eZ�0-�MӉ�%��R��<��G��Mx��4��+��S�d��d�Bt6�LfQf�<J�����a�I��j/�b��#��U�p��ښ� H;�2��^d���-�H�2��4�$�m_���2Ne>���?`����q�TX�����1hDH�U�tNs�v�J�sH�,``�i�x�]Wu���MKY������.%�2��T	w�%��n��[���=���xlm��b���PFCL\�ݕ�:�C��#�YP֡)x�� ���ODN�g��?_=��󭮣��7󂈠=U��,i~I��'�a8�Hl_�����r��>�j7^
������,DfT;��uH���w6l���傈���P>m�,h�i�+��;
#��c~x:t�p�Z��������*;G�;��&L&�ҕ��唧_5�'/\��VN��W��wz���a���@a�����J��'�yk�R�ba�j�p�s<!d��N����X�N����]�x�$'���I,R��'���>��vS�u�,N7���KPж Vv���p��(�|�.��ycj�*[�#�����:�5�O8b��Jég����61J��x߂*@�O�ga�4
�2e�x̲���b$�B�������qtH�g.y�_��uV��^~s�]�ʎ�<0�)S4!o0�G�k������	��%!
�o�&OQÿȸZˉ�.��L�1�1��%���$2[����ADPs{��tب�^K�����0ӹ�+����Ԃ0wq��o�\�1�x�E���8�3�Z�J�WB�O%�O���|��<0�Ȕ`"i��(U�Z7oki9y�~l��\��,�1�l�!i��M�m���\:�ps�) 0M�$��lw ��b"��3��B�٦E����Xn��"��/��|�S�.��:�v��.��ے9�q�ŋ�:m��%{R �jT�H��IDO��ւ�����u�n����>(sx,i�CR���V���{�˫�\�R�fQ<[���>�98��K�KwXa�ݺ�1��X�p�gZ���t�O���$����VuX��eC[�]���f�'T��<�Ik��{��dF��B���븴��)aKTf��F˕t�<;�i������eo	�(�G��E��m�ϒ���{+��q�f?���`���",r�y�y)<j3�7a�J϶�"�O��x���t�	G�--���1*�F7J;�nO�&k��'��ӌ�v `(�
�ca��יgazom	�C�B?hY:�X���M���)��$���w�jk�1x��	��ψR����Ts!�Eu�wv�� ��=y����v̟�H3�fMP�#NK1�V`u��*�´<�7صm��Acڬ ����:'r{�fH��ڄIӰu67��a��w��N���I7@��ˑ����v���bL�3t?{��=��D^�-���[���ͰKO}�
=��kuB3*�&���
7Uz�?$� �ys���t���QI9�B�ڷjqג�f��D�Ou1��|Z��U����$�0K����g,�Z��h�M-�^�j�j�ޟ��.�d+�K�2�L��~��V���E�H�{=��iC�ځ]
���,R��~dbB�)? x9@=�^~g.�\�X����╍g	���F��0��}JHM��X&͋��g!��E�v����Ax�����xIB!�پE`d��]f+O�
�j�!�c+�Ov�q��3��:V�y�f�	c�w4��#Cs��D�Kg�(1��x�f��A���ֿ���U������W!�/��Uʈ�MT��r���2�P+)ִƓ'Q��;���&O�����do]��Q2$Os�pi��M�Q�3��E5�y����\��%�?��)�~N�=α�9	��v`z�F��3�mө���Z8<�>��/��������V�tIP,2զ��5��6Mo2ϴ(D��B��~����ό�s��`�jon�Q|N导���+�g�&3� b��o�@�^�/�X>`���MK�>�� Ia�v\��\��e�g�4/�N���X.lc�ٽ9Y��a��:�:������Pq��Q	0�oJ՟�׫Y��w���Mo,Sϩ<�d"u^x����޶�H<�ׁ��H�D�f�s���x:����|�ư�)R�ےq�PH����~Ԏ���l��QC�_x��r��P��;n�����J8���\����v���Gs$#k�'��?��K�gS�gw�Hl�h�FQ�!@|��r�IA+k��oTp�Zi4H��7�-$(^��m���_���G��i%Ɂ�m�v3%��P�2"�!_؞�^Z �tpF|���N֩�'�TC!cP�ο�;O��O����Mt��5�:�=������Z�BD��G�0C�]K�(=O%���ns^�G`����	H�1kjB��8.�9߭+�v6
;J0�'.����W�5;�z��8�)���}�����Bu�Ή�Qh�d��!����~�����@G՜�O���b�f�׶����V�GO���1-+ffc$N�ջ��l�52��E��P�y(E3�����~�l��W���앐�SK�c�������2SsAۅ�\�K4�P���&L�4�y�9 c�p���)�'��2V��2���;ψC^
3�;�r:'��cM���M�Q��$��cWT�9��n�1�\��8�h�_w�'m�_� {�}�R�ނ�D���~�5�$]̓M�'� c*��-�j�P�:һ��Q=�͛,ꆉb��|L�1�H�=W����
Ra����Y��NI�n�t5����Ż���Đ�Ho�#��O�3�O�,Ꙇ�jex '$YS����2{%'��$�.�_����V��BH���N��SūɎl�^(��c�;"��Z���.b.�"o��?�$�'�"!ǽ��?����-��$w�,&�γ/jh�I�'��� �Q0�p��
��/Z5�J��J���Du��*��N��S���^[0󯞑�hvтE��+���LL�Ԡ�2���:�����%A��P��?�\ju�rqP�}���&�%�r]�}�P���Bb=�m�J�ju\��ۿc�$1���p�2G	�F]�4W7��?�^���g��k�3�SDhP�um�"�blx�,�ِ���v���`B�gB<BLF�\�fw�i���Y���������xa����a�sb�8�����b@"z�Q�?&���t�P���*[�\�shԂ���HҡX�h���p��	����`����T�ȫ��b�Y=�������v���LоL~��U�t�dS�C m��6� �EZ`���Qlo\�&)� m��~�dH+:��܀N��Apc�g�V 	�4�-_�я�a ���&�Aw��n�!��aW����%E7��(7�J�˭" �i��:��g{�.���#Nv@Tؔ��j���=bz�ai�!��ط�h� ЍuS�Q��C+o�M���Ǚ��bu��y��Cf�պ�,�Ĝ'{afO&�2��@�H��ڀy.Dy\��O�6�����D0��.�Z���dK��`}^9أۛ�{7���3b���	���J�u��s(��	��7i��zIɪ+�%�֟Rr�����.DO�$6t��,Dy�:�_�rfQ�ī?����1���I���f=�yߠ�<YT��%�@Vms!.P�L�=@��8���~m�=%њOf�\�c��j��K�ߏ�63����8��THXdĝ99Fg�$�|֨�JZ%�v�\*���'Ԋ�,���VK��HE������ng����ŉ�d����1>���Li*6Lroc����χ��/�E��E7�ϳ&�]����'�I��!�)
]���2iܣ-ˈw��\�`�.z9�ҍ Zb�UN%gz�@� %e:��w�3�,�ﲿ���oKN��e�5�,��9v�I#).(��(���BʜL�U���*�ᇧL8HO��H'륱�b�"�d�϶Cq�n�Dv�5�ɭC%�:.�?L�És���݀RR<�(S��>�T��r܅}�#h`mgIJ����F}b��©���.�d���;P�m{�"����pTs	Y�����h���a_?�V�o#��s�١E�z��p
�������g㖥�=�-2�����me�%��\��Rė
�/^ӟ7�шgL:r���4"S*u�r(Q��4.
�믆�j���6�v�ΐ���ᗣO�p{�l�꒎�wv�Ӗ�+ҹ��I�S��4����S?U�� �g�tK����I����\>9�#����s��1Kc��`.S#�9�D��ǞPAW/��чfGE!��R�
��'E`� ;C�s(�c��mY���+�Qw�<�~]��*���9��r+��,�����X�ӄ�٤P]k���	�6Ezo�&�0ע5_U��+�c���8���X���}�0�*��z�z"��\'P�}�Qge�e�
Vk����Ìw(o�c/0*s�e�?��x�X�j=��f�z��^I�����Dr��*��+�T��� �CA?

�O_o��&�E e�uhrTv�lP��+*�� ���96��ē�f�M����]^�F�_�T^�����`�(y�
�P�&�?�� �Rp�ꦡ��K�����q:�W�THN�>��R�Qr���R��]�~P�bY�ߎ������)���q�W���fhW20$	�φ�)jf��
@fK��&ͤ̀�TE4��W�!���֭��y'섄��v�H�3i@-i�^*��e�:�[�4,���5��Yzy�'��>���MDeO�k{L���~:���
_�R��P=��R�nI�\r����v��/]�q�mey2��q�.)�	lkV�8b,|�/�ʫ��W��;T7
>���Df]���h� �ǹ�x�xP�6�q��ֲ:͝פ�`J����d#�'%���lgߗ�,�?ҷnrN���9�k�WV�,�i7-�]���:��&J� (l�����
O��<�D��ƮVl3�c@��p��Z��}��;�qw�˝��-�ҍ|gF���׾j������O�U�����!&G}m�'�Z%��n�G�72IY�����_�i�7��%R����%�(e����=�wj���'Dؚ�8�@{sh�����E~\��,A�f��;r�V(������+%��Q�ժ��"'�X��ọ\w�$͞��}��}F�����5���:� m9T�?����e���^��g��x�5�;�Yɳ*$��k�*��T�cd��juP�s�����G��7�L�x9�I�#���;Vh�x�"Tt �g�=4�2��U�uSc���B�XkQ����������ӫ�����gט��P�Aoՠ��۾�>�j+�R����I��i�n�P$�.�������U�%��Us���]�<*e����]�	�'����'�F6f�����.r�ڏ��w��][ �����}%������,��#�^��'+-;�VA%�K�]M�`��.LY{��t��P�z2A�i)}NzoM�df��?�����b�G�q�O�T�I"�8���jn���7(�(<�=ᲢO����:˺V�|�o2�����Ԑ{�f&��(����0*a��������pw�<J]u�ls�.Ğɍ�
dO�&)N��؝�W�'�]��H�ouʟ�c�[j�Uť�:G�3^�ؿ�7i���?Etp��W�_���,ؠ/@a9�Q�Q��q��w���-]��"�g���㣊��=����M����7����K��ǂG�X�G��4n��wډ���Oz����Fخ̕4���`5CD�(��X*P
i�5�ߑ�?��`4 tM�3�'t�����k�Z�*��E ����\�#%�E�Jh�;)@\�ǆ�0�J��( rt��8^�K:���|HK\!v�ޓE%k|�59�x�,X�vڞ�e�q�j���v�"O�O�����!3����m��������
�kX�/ۭ*~L7��=)��_��?�ʒX��gv��yE��O������Gf t��C5��6e5����٥%�:97���7�(�d�T��Jƈe�;�qu{��m˓�c���1�/0��K Q&�cbeO៼��� e%x�W�S�om&2�I�Rm���Q[*�lG=ߝ���w�~n�ݔ�l>�t�sG�̖CW��1eő/�-v�ʦ�(D�Y��C�1���U��!�Ӽ���$��ō��C>	m7�ߠ)�>Vy��g*2��G��]����&�7G��D[�r������^��[D;�sWf���eFv:*_���x��.�a��3�́y"��_Qi\|	g���Z��}bt��)��P��᥏d*���|����`w+a�ѕc�AɌ����t�!��*�t��@+`YA/�mhy4�*`H�߯}����NA��<Z�gP5aR�=���T���Q:�!�1`�W�8�$��Fϩ���􈏇���K�����/ۅ�vՔ@�A�O�M�(�÷^�?�mf�� �{g���$�������Y�=��‴z\�T��[����FX����F��������Mx �MBĮ����?�+C �a��]}O�l�#���F(��
�CH���HΏ�K�F��[j_��?�!K��L���2���܉�k���.>$}�u;d{?F��������[X'���ˡR,HeS�&�T.�*�25�gMv�_�8e|k��+9����
c���y�Y�ݱ�媾��é ��E�m[��d���XjГ�~b�-7c77P����.��F6A����ѧ�'��C��'�3&jԸ��r���a�'YKʐ0���2��>���,I�j6A�N��X˻U��U�`�b3	~��)a�'��[0���'��1(3����8'D��p�J%8���!����?^ːZ��Qb�����?�%��]T�k�h�6YO������>���"*������$�Q��?�<���|`$�mJ�3�m��#1{_����1x��c �qN3ܺФ�ٮI��r��kRY�'T��a@EM"t�\-	_�U�Z���3�r)�ѳ���!�=�ԕ�����%�Ē�b�s�Y���q)��ʅ'M�ٶ�T.��B�V�?(���O�eݿ6j�ڋG�öV�)���Y��7]��Ϩ�oo�>�B��y�v�E��H�+|/08?j�u�qQ��7Z�B����bjW#`P*���)ߧ	H�H7�)�)��w���;�H��7���܅,���0JPDltT�'b�9a溷޼i��K]���#��P�Ӻ�I�9�����t���B�U�0�	x���s��}�:>����4�e�a������r3�3*��&upWق?�n�	�'F����4��T5�0����Sj����(\hM�g�����9ք�V&����Q�����HryI@,��2��7vB,?���b�r>A�� ����7�N��sC{�ß����m t�k�-����xy�R�V�"�#8q��*�Q�l��U�1k���\��Z)g��2]ZK��l��8�C���fs����7�)0�b+N��#z�Љ���v��h������)[N����̧��ڐ���zs��3�i�rբ�E���{�9�5v���������F_�tgXR{j�d�6��%e����|M���.i&i�7��\Hz��̶�%� ��Z�_���@��Qdz�c��k.��[�;N'ΐi퀼�r�\	�t�S�9��y���p]T#6�Ⱥ����$�ZT�$,����~`Ι��͂'cW�td�L��\m�zɚ�/��Bn?×�\cAP�Wۏ��[����x$���'ѹ�@1��ǿ!r�?�D+\��R������O5}�p8zlz�QGl'p���(;U&�mD@S����~�Z��h�=(^d�c#��bځ[�Ό=�|��qF�C�>8f�z�+t�S0Y]�0�`�ݲ����!45+;�T
��`s��sS��
M��B�W�O���9�܆��pW÷�KkI�oY�]��u�kp洈=���L�lE��-��4Z�&�o�Ru-vO����a`A��^�����q�¸')П���1�S��lp��|�?�pǀ��A�'�js%n4�hȷy�bF�u�̤"�*J�htut��1eN#�^�pX,��"7�Jv�\�5���O#�K�1P4��hB�poho{������tѱ��Ҫ�6��6������¶������	��ϓ���D6��K��qr2|���i��]WFiT�~���RrJ�V��0�B	d��O
�i+�_%�6���.fP�ᖪ8#��:L"�qi�YMP�H9@zR�)#��.�-�L<V���~e��@A��F}��������;�'�(��h�0������(���feeҟt
�0�.	��v@e�=��!��<qi��:���^g�sB	K����@Jy(ۆ��]��Q_<�X��.�蟕T���5����P����N���3�Q���1��`�c���*���|�rtc3%�W��nTCJ�ޕt�#��P��6ߗ�R
��J�#J7g�B�>�f�SE����G�z��YH�@���'�X��tćXO0#$B��Y �����5eJ��
j�+12u�-��cp������b.�*go�_��	�ܝ�Q�"����DY
����=V��^0����ٰ��2D��2�~E����W����Mum�h�,1;�l�4Rݺ�rĦM���I���x���]Sɫ #6�d����j�C׋._0b���������L-�R��u�E¸��~��.,�3���sj(U#��Jz�a�׎�+8I��q�?$gZO��
���n�1b{��b�U�	��l�a��syvy�F��Y�2Cw�Q�b��lz�b��j�#2H���	
"!�n�<� E��N����+k	̂zd�چg�T2���^���w��kVpq�H�Gi���,~�,��J����ʒ*���5��S���jn�BAT�i���]�~ҍ�R^⍒�u�\
xg�<�#�Ҡ���ÖA��E �����rc�{6��"� ��"џT��>K�1kx�������XO�:A�H�G���a�ה�hR�f=}��$7���l�� ڙǠDV��`���+Tq��<�H@`66Υ]
���e�]��#<ɤt<M��]l�^af�ݾ�u���_<By<7�{���2$go�#a5���J<��n���k�9+1�o0A/*��'o�T�D����Y�����Gf$^U�骸:@�����"�pO}+큌m�~�6|l��B�s�PA��z�9��uP$�G+-@�Y�t�S���'ߺ>ݘ�R���+4�6���B�~�<��>W����D4�3l�� �:ʬ������:g��i�;����p����2�'��_��ش��-��.�A���oĳ&uL�y겹��xSs���b=¼~�ek�`�nu�n[�2"pӃ�B���>Pkz}NfϝZ��(=?�bKv8��1����FM�p�~Gaߖ8 �㳘̓]�@�w��W�����eΨ����fe7i�	�nSx1*a��p)�G��6h��z�.6�_S�ͱZf���C}��l1m�,-g~��ax1������N�u�ப�_tJ�&� w�\j{DDG)_�`Ǝr���]���5��WߐV����E�db!-r�V0��d���_��0�pu0!ڢ G��&��8�L#[iq���0�����
e�|�uT�Qol#*Z���o��W:N���`M���,�I���s�߇�>� ד�%f#��6�7�'�T	eö�]�{�W1v!��(�l�~�k���T��S'v�������) ���m,�9`�4:2�AD��P�4�ІՂ|���-���rÝgj�#�Z=�YW`��E#k��H-`�B�\�)��O�1�Ng�O#0O�w������
�[��'r{���ʆ�V�T};O1t�y+�9o��-\Kz{���
~�&�����7�;��fc[�[��{3A��E�Hb�1b���:�fGI1bO�gX%8�����82R\���˕N�؄�e���0��ߵ���k��^�oݹm�nTRGl�櫪�	ѡ�V�]E�7]�We�>ǖ����b^B�� �yœC=�+����_�,�~��!� ���66�h�`�`R�*�^'_:B�%��1�3�ʛO���EO�j♐ۭvG����_I��>�:^�ˊ�2�����Fa�o^F|�I/)r�F��fȶ���q�J��ب���|�������+2T)��id^X�>:e����n@YnF3V��Y�"(�ʹ����p�UlQ������7�����H(2Y�DU�f��A�ʰp#���J���zfU'���r%�0y3�,�x��qd����^�E������t���F�P��گ|�Ĳ�5g�,D D�����=�W�ѕ	f�s�p�C��D��m6D��P�b�j�A��������t�޵D�-fK4>�^nZ��UG R�d7^^���v�
p�|K:?�qa����%l�=����f9ƯBn�޲�_n{�A&H7�<r�S����n�F�t����������nO\�TT�C_;�I�
a(;�S��j]�ñ�^�u����Q�������6��8���¾�=���e@�wb{z����^�oh�~�(q�f��ԧdU���U)�֎g�`��LV���Щ��d���'����)��9��Q%�H'=�BP�&#u�K��n������<����w.L�T2�'��3h'�����:��Q3��|�;/_x��r<zo��zh�]vQ׿,��'cU$���]��ۼ)u��$}x
 ��m���p�=̾U>�l�x��YL=^���^�\�S�r$�j�^�SB�2"bmr�6;�0uvҭL���"�d�@��2b2��)����OG
2'9�O�+�X�p9W���cl����4�d����쮕^�� ��"Ş�+�4={�F?�k���١J�������@�4�1�E���Pu��w�}�� �A�����ْ�I"z�q]��a)!7�&20����tpG�:�39L��z���B|A�g*�=[DJz�f�i�&k`b�xս8�.ĝa�q��ɯÇ@i���ψ^^MO��"�����Z/�������#Z�4{I����@��i_ecє�D�m��)!;,]U��x���k����83�Y�֑m����x�Nj��O�]��x�K��f@'w#;�8��"���&�{׍�-�0�J?��WV5/�%�DuM�M�����Ԍ��G��$�p�V��1� _@�`[��'���(��j��m}u�!�@8b���bI�����{�I��=aQs�Q��>6ct����c`اR����O=B�A�I���F�-^�C�V�Lk�o)��NBJK&}���c� S���1�:-H�o�r W�N��@]k�rR��SQ��G�{s���\5͗4������E��膚'�E�{��\���xV� �^m@�#��ƼX���wF�� ;���[0&�HxG-n
%�����yƒ!7�5��\$��#y�s�՝�*�����
O�_��O��v�ԫU�DDT�� ��^���YAY�����ʞ�1�]�^��-&�	 ��9����i$nL�h����߿՗�Hq�r �^X���rVl�8�G�.���!eD|>.���ӍE�{B�(0Ϥ�o��hX8N��G�Y�^�N������bn�|m�=EED#�T�g�Ǝ/$�b��۹3JǮl�)�[�9�����pt�5*:�������K(�~���3�R�]���ˍ9\�=D�#��h�1�� `����?0pa����j�������v]gIo��Hrs�.����>�7�n��?�~��29�?=8��s�-�{PD&�i���S�?~��h���BZ�8�����o���Xق��Y����[��Y8L��`�+*�SI�<����cW�?(!8x�E�>�%c�����Mw�!��zʱE;���i�-Cc����xZ��iq���n�b��	Q�����!Ph�%([�����5z�ё��3o��C�'�{c��x�/�G Ї��9�� ʦ�����F�4��-R�!Ꙑ�d�h�O*��n��x;�_�sȵ�W=sH���;*B6ΐ��+s.n6��L�$�C"K�p�����,-\�%����B]�K_|�G�a&`���g)@�s���+��Ǿ�t����c��B[TGZ�T�`�� +���aC���\�U9"�^����g[e�	gŬs (�f��6B!�!U���)�W�=��G��^�n��H���(�i �g������_��#,5��$�1�^�C�v�y�PI?��^�s�Д����Z���Mf�ܝ�:��ñ�?���^�q9���#V��y�櫂�α;��?��V.��1ŕ �L��ӸV-���z�Qlb]����	���=z2�Z�a2�<i��J�n��t槢~ya�؞X�z���%�'�X`>C�}�O����=m_!��<��un�R٬[�����e�āw��; ��ا����zZJq��ï�]"�J;�	�Χi�!��g�)M&��_K���g~�<�����G�����>�8��6��� ������ڄ����n�� ��Y	A�T��d���T�K�ܼ5���P�_ǀU�,�6(yɌ!����(֛[�	8�+X/�u�4��.�W:��R��ԵO{�m+|i l��N�?�g������d��'��vm� �u]|�Mg�[�~����/��pg�8
u���Tt́X�|)xG���&�[�h�
�<�|��8ɠd(M=b���SU�)����f֐mX�\u���\�#�ܧ;̝ �C����BvL���Z���,�R�C�V�=���op�	f����s�/7��m��C�����V��W͘��BK1���d8*?ס�$e�i�>�������1�a�<����aP�w�T��ӔS~��G����""�Eզ�������s�������:�i��*����)��	��F��^���������P��Z��--H��������ᰝ\�)@��#�|�C^���*�U!*�d��[d�"(c'x��F �%)�4(���,�BZ�w��o��ZFU.l�&	_"���ҟ��=�%R8N��7�	���xNo��-�D(O�j2�u �25~�� �Kcw'�LX�^u3M5�k��&6"�w�,8z3G�P�K��q�~�q�a�Jd�g12V�P�gJF�ͣZ^�&M����k�j�Z( n�"���{���A�*�>��\l�*�=�ߞ��1{)R�]���9�W��]��{t��?�3��&F>{?Q���?%*�x�k�Sx�x�r��zErz�@2M�Tހ/�1	Ra�	3a2$ 9��H���:~X-ыܘ=/o`�V^�-��Lk��=f�� �}��i땮�蔓/�F����hY	/�����ouP��f('�?+[��͞b*�$�-���A���؆�
3���'D��̴ ���uo�?X�x����\�jHi�aP���J��E��w�L�4GV����H����釻Y~�02 ]�<�0�k�|�s+Nx�\F�F�d��/���v4Â�'��5�5w}�	8t�P��g�uD���D��s��;�E��ھ��ɏ�>��+d��B�3yP����������Cz\�6X���e�^Bj�Vs^z��P������0�(�q����7H+�w�!�W�2JL�D�O�����.�c�����,��q`��ƭ%�%�\e�EMJ|Ǳ��@�'�8�S�z_�������J	�Q=}��ÜF���*&�G�-H�����sf�!&�iJ��(57Snm�~h�lq�m�EW���^����h4�In��<<*�{�D�Q�G��'�d?\n(�9CH-�σ<E�?{x�T|gF��o�~ҀfHϤNƷ�r[\6���s���y5�O������L�>��Oó�>-}$wRy�[��ks��!���po�����N���� Ӕ�'/������p6��.l @`��S4#!6��קNݦ�:�~��&����o�T
duF0Me`u�'��q�!Y��6	�B�lpcv�\��'H��Dj�⢙�G�aM�n$���{"~o��\&G�mg��9p���-{jҿs0�=AF�y���x��rO�SD�d]��������}�/ʹI?0?�C� =�*����\���h�V��Ӈ:�aYp�a�BX
�aw��'sE���$5]Z����E��(���.d���&��%�wI�#���9+���@.yfʔF �ܛ¡�0�u������^�e�@�Mufq�ƥJlg��؎�H�"��e��b5-�̇��.Wa���Gfכ^�U�W���@Y�h�����g r�$QW�	@w��B������MԪ��aE]�_^E��c��P��W�������>���䕶�c�;�W�@14�ˇ˚�6�[�At��y��&�g�"�v�)��U�$Z�y+����G��
��d�ZC�\�y(�-uƉm���	f��5Y��� ��>59���O+*�����嵭Qq���j �.g�_3g�[Ui�����\�p�@��\#ܔ���t{Ċ��2h��l/�e��zZ�y���Dߴ �}�n?��X*_��2��xl��K��Ę���[��~����:`Z�nz��Ğ��jl�'���:�T6ծ�����qT8��b|cw+XǸa���#R;
ַ�����]�1w�IM|�f�<}#�n����n��R����0���:D�C�.E�>][l6��{�ld��5Б�<r+Tp�����Z��Z�7���f�P^Y�'�W1�٥� �(Ӡ.#���� G�"�jβǯl�!0N��"��������������T+�bj#��D�7��ǻ5p���`d��/�I���]�(�Ѩ*E�+�2:�U��$K�R�Q(DY�9�?�l�+|h���� ����3rK���f`9`�f������}����G�y�˄����:�����RV�B	�t�p\�����0�V�0�v�ⴾK�y��� /�o��H"��)�^'b� CJ$�hʛ�vFv� .���6bf�,�ܳ�0<�:�V&q���><� � �WS��ռ"�݈�r�F�Q7������
Bط|  <�uK��kN)��� � �{]E�(�I��kځ�˚��fU�Mo������	�R�]�tP�����)��$�y5R�=�t��0�C�zNn,��+�&Ob1�y�Q߰G�/f>Vk��>��c|�u��:��0E�S�_�4R�����tU\�_��5��1{��%���c͐c!%<���
[���N�?���+�陋��N�rZ��6h�f؈�s�\���\='.����5ANtP;��A?���<ȍ���ې.'l�y�ǫ�in���# t�ʄ4j�Bꋞ�!f�3�;��+�eARP��r-����g)�-�O�)���%���j����~��~��=l��;�Vc��`���	�@Z��KH���?�\��f�3*�wq��Q&��-�� �$)����J�w
e�}L���-���D���a�@k/�|���4��K���Y�[�������*x%/�ȅ�=�;��6�W5��ж$$Aj|o��f������y;� J�C�m��l�X�}D��Z+dO��mlul%I�q�=���m1Mp�Q���ӾT���Ү�T�g�GN[Ck�xH�yT��͘�\�.�G��^�R=<KG]Ms�m"��=��������I�c�{�y<bw�7�����fa�xఛBƯv���8T^@WՍ��-���Ѵl��2�H;�N�/�pSG}���4�8�[\�{��i��	a5�S�]'��u�b�yT�Ν��A���T�P�kF�dt��Q�	�F�iL�}✲į�/ƈ�k;�25})�WR�7�֥�m������9��P8�GaU���)�����	���z[�~Bd~��~��2%`�XAUѵ�bQ�tL1� �r��J�s�6W}�qn&�����r��,Fe�틮u��&��J��=�Y��:(�8@o[���q���7�P����s�:R;i�oˉ��e�B����SQ^G|�08��X�H�F�,G$��_3/��Zt�A��h/���4��#s@���k�we�����z	�����p�kl��3�m8�R�s�"s���D1oj{F�s?��e��w	 ��h�|�����[��`n}�F%YUU�QګL�S�Г��
Y�c$�G����eTޅ]����{Uw�C�弌2J�$��h�$�����sϕq�f���I�L}��AJč��C�:�j�ԴD%�»/�$��c�E�~	�s`����
�c��$���9��{w��N
�������"��jɐL�����q�O�q��Axᴜ��%D�S?Y���H������6,v�z[�������YF-�"���ٝu�k�x���/�ft��?�~#L�D��[�t�W /��-]z�?[��U>�5�	h/~o�P+��t��2�.�	}%��,����9�=<�h�����MMGߎ��f�m��?#�S�X΂����#j�$5�b8����1"wX�i	DJqcMl����B�WKx�7�8˺2a���of�?��C��-���#T=���M#S8 �����A)�V�;��IU�s��H!�g���$�� &�c{������ҝ{[�_��i4��%�s0�L�O�2�A�7��Ty7�
����K���p��}K�¥�B ��t�9��M�;���r~��O��W�vꍴe�LȇC��m��tM����ZI�[�=�o�����-��ܤ��nԒJEsm��P��������1s
TP�A��dH����R�7LS{ll!�+>�ӑ*�,���p��i;�W�E����0��{�]�꼖N �V��Q��I��>*�����2���`�;�G�nj�#�y�:&�M��5�~[\ٽ��@D�l��m�9c���J��[P� �#x�f1��˲�N����¾A�1?�0M���[�S���$��?"v�$ ^�I��C�-��D5�K�(y�܄�F�a����Pl���3�~.úؕTwܻXȃ�G`SГ<�"��®�|R^�zKY�y�w���v�[1�J.����f��%�z�F*�J����L�B���B3���dp��,I`D�+^ħR��ŵ3���x̳�b�@Z�طD#�{P�h�mcD6��	Ѓ��g�}��GCI����h�w�G��s�$R�k��/K�7���aV��h����7f����n
t#�PYZ��$�E�v0�G�y՛.���!��$R-�������}E:ߑj�8������6&��|���m��
�
�2��M�L��u$ʖ˭�fY�f���Q/ʠ���Y�3����&�Ʈ(�U�_)7ۄH�#J���=��5ϓ����j[�oѤN�p`1�E�fd������R*��B[�Sv��K�-&����k{]�k5:˛��}������� t"�oq�3�T����H�q|�>�%:*(#��fԄ��͂�g�Mr��2��.궞ˇ �F�/�)g���q����4M�Z�
=`��x�ȃ0t<g�I���?y�ˎ�h:����ZN��n)������h����w���APx�F,1������*�@���t�zh�XR�ث�a=�w<��"iP�s.�^�u���p�+C^�B|^f3��5�ssj�5"-�/�7�������6��:he�M�N�m�s:5rz�E1�8|���|ɲ���w�"����LP8������̻q����(~X0�}ʼ��	���,r���i�ۨ�EԖm���b:|z�P1��o��M��j���J�JP{�Z������� �랋.���gq<e;ݏ���B��E��Y��G8�Q���2�'�a¤�b98�����GvR���k����m��!<zE��� `����m�n��!��@�/lb ����E�V�]����W���%%[}~sa9�-�~�d�����N��]��*I�5JU�p/��e��#3�Ķ-�d��m�+�ښ�y]��Y$L?�4��;]�xޑ�fS�v_���?�������S��|�]E.�2�܇�6Y��v2^��ewdX�N�x̕R��JM�a��^��V,ѽ2��oq:<��Q�qC�����5N�|"O�/ڃ��=X0v�N; ����0@)Ɏ�ق��'�n�Ld���Qs<�9��)��8&�= ����~8��5��p1�tA`]����4���ϗ<ŷ��ڟ��sE9�p��+�kK��'��C�W[��8����9M<@��#�#�{j�$ݵ=D��V�L"�R�Ѐ��	��vN�k$�zުQ��G/�Y�!$O k@�r�Bo�c(}��w��t�y.����	��h��ur�tN�� ��@�W�z���*t'!I_��ϟ��J�$xƞ-i���G��/.R����'������3�)rm��֟
g�m��q�khg��.Gmc��TF����̃u�K�j��bY�y5��{H�ƛRui��V����6.�lݩ�rM�_^���:�ծ��p<74D����N�]��dqT���"�������7�?D����'��n>R2��?��1�4�Vx����$�Lh�B���OЪ�Hg�Kk�Pç5�X)����д��q3�z���� 	Nf;�K���8�;Q�G\��2е��>.7�p.�57^��$�4ǋ��\��_R�闸��]��ߋ��~H;�s����wD�a�U+m*J��"9���V��jGj���1��1@u��	U
�\�	��;O*�C^5/�H��SOM��{H�����B��4�5ӓR�Ufe��u�k��7�,#�����j���bI����0ya{v�0I�ݷ|�d��P�JPjS�_��ޯ���Vۉ�a��L�3*��*g!�� _�P�����U�*NoWE���32׀�::X������3�<�QH����ʏ�K,�Qbi2���k/��BhPf$R�[T�+	��d�D��	F<.�I��@�&=W���i��`yȘ&0��͌2r(�V~P4�lO���z�I���@1>�ʫN�>}�'g���^�! ��4�ꂋ-	�ɴ��D���