��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&������*��q5Ji�6�A�+�Ak�ŗ��Z�h_��f	}�G�@����Ԟ�������f
��kRN�������pm�bGCA:T������Z��ޗ9�Kl�
�f�ⴷ�����s�`�@����X4( ^v�UWP;���;75�U�
�\g�vC�HDM�&����H�i'�������>�M����n2fч$42>레Xɲ{�7�86޽��/
F�eQ.�~��O�rꢓg���@���!���@�:m?-T�{/����=�y7j!��#)_��A,gS{�G��,�1qo5աfK�b���БOJy4��&���\�Mǂ�zH��l>�`�J�.*�@SA��-��p���>��]ήq��,@�5vzV�����751����3���]��o��ڇ�P��D�d��l��t�3I"X�u,N"Z3���ҽ��N�¦g#I�EAR�>�!�O�cl{:�Р�Wtx��5�$�9���&Ha��(�F�ajk�#�:���c�,��f�A��,m�6�F�]%ү��M.0�%[Q~��A@y1=�����3p?��:
ʆS>W�wC>�vD�J`o�h�������|20t�˥����8G�{m+���m����R�M�:�葋�W� �E4�c�>���K���nHY���'��?Vщ�"p/�ysm�;7���l��
���&�W\T���y�E��w�S�>#��G�R�A�)i����5��CsP�0/�)��M�ּBO�D+]MW~V<��h�7/qZ^DqB���_��?��t�5��;��G���:�y����9)����������!b��ّ~]r"�j6���aA6�T�����R�8.����O)�Ļ��0���-TE��I�l��T�<��Ʀ(�G�&��	��L"�R�J�1���S��<�YrZ�K�q�l8�8TJ�e}�EbLZ�?M�[���j����92�rd�͏�n��z&Br��mV3���g��=��@�𦈇$^_'�8��e!4�g*��Z��8�5�KܢYJ�o����&��+[\=n���g��1u�0��=�1M͓FC�R�qz9Ƣ�)��i5诵���}|���C�J��CTWl#kFM��潋te�
_Y��!U%����Ğ�go�J�1�ңx�o��&jĽx!�������ɮ;f�:�M�tFF�I�?�\˜'�ɥɠ����;��ᶉ\9:�9��&U�y�W<�7���g�}}u����y�[h=b�-Tɍ�ND��kVg�7�@Jm��
�lk��C�4�8ÛVntY���yk���i� �)w�Ó����2��t�%Յ@��s�B/�/��G(��(I/�C� /���D$��o�S���
'�Oy��,*Hy{��і?�;,��h�����ͤ�O�z$��yqa;��}�|]��4*��X?#�]�%��o'��e�F�f����}��� �˞���N�G��{vOdf"Qe��w%��,�-�"t���-�e��9ä��wa-c�Sy2JQ�
�:e�n����Rx�#���qڧ��\��?Q4^��W��QZVq߭�O�G�?ᨨ��DAhcA��|j����^�:��X�B��(JY���Wn�-y/L���k��)������ϥE���~����`���T"�FJ9� c��1
�pI0!�.�|ZXeޔ �"� ��.!�m`�Q�Y�{Ri�?��h&��ǁm�Iզj�ˮ�uUlB?}w�j�����!�����R~�V��O(�v0�F�����	�R���ޅ���Wd��N�G��
 ��Mn��"�mȿU�������>��l/ӶSg�l���#�4��>}`1�I�F���V��;�iC�n���j�~Z�A�&�]���^ʫUݜ-��AlOӕ�6�32f�wo�f ���H���i�o	ߌ��*�U9��q|-Ɏ-�(�p�/˦2"���ࣦ�c6UyB�n/!`�^�_~��	[��D^�����3�@����u��{|ux6��KÍt�;��
}�w) $�������hY@ m_�]����^-���	�q���3����oy�m�)���A���GJ)��?Mo�u<&@֝F�+���#���6��O$���M%����<
P���̖ѭ˅E����O;h�4��VM�a5�"�=ts�2��*�g�=�;�K�je�̝���0��Z��:e2Z�� %�D�I�7�*R��k��!i��ϰ�Ԑ���C�6�J���cGŁ`3�\h�0z>���ˬ��2��t\��:<omfǥy��|�}V����`�;<+_Cc�ʁ�,ǆkE��{��d(�q�+T�݀2^{9�����m����_Q*5���{��1
 ӻ��^�:_��{&�U����:����#r�U�"^�*�Έg�[�c����C�$��&���4<��dD�G!?!���K�At���_'�:�t�R���V; Sd���1�SQS���>�&3�cJ��9�����[兎�a*KU;f��i`�3�
C�]�Z��_@*�\�$�ْ�v��J�r��@4ל-�p��0���]i�RH�6Au���R��(�j�V^9�)��3^'/��)�>�na�c���/?�U�\OaQ���U1�ܻڤ{�	~�x�b��R���+8Ҭ��^���qx�d���Qړ���Q��Z�n,�2�8�mS������)-)p�a�
�EY�� �֪�2���X��7�>\0Sr�����l�~st������ǯ�3Ҫ�@�:�����6�c��=����MO��?س�sZU% �y���1̉�}�E����\��cZ����dg*"��A�2��
�(1ː�\u���)DԷ���s��;?A����_E���� v�(Q6� ���LM��
�O^
�ͱ�4�I��`� �D�T�$%�Q�]���F]I?B힟�-Rj�J�Yɂ?h�@���¼z~-��&(�/O�>�ٔS�$ˈ��H�����Sw�c�P�f�N���/�ڠ��x2���_�;���c��b
 ==1�tܘ#-�*��6bθ�Z�4K��O��Һ@"�8ѧ�_u.���(y������ �5 ��p_�.���-9-�׹v�fn.C�F�fZ��Q�S�[��<�"�X5o�^j��Hmv�G{�֡��8�E;��1��`���{��]�����Ԋ g��z6J�3��
m%�uh[T7�%s���$Ķn�os��k�+���kS�p�j	��#���u�s1'��gU'�1G�3���o���V�ֻh=KkWK������lE��aDU��:�n2�y�*�/Hj"��6��DG6+�x�=Z��B�0/R����AVz���xs����)N\ε�w�8�/�ۗB�ޕ�/�*���V{I���E���Bw�����4��6Ri���"\ɸD�eOr�8j��o�W|�r٣mr��Z�]��D$ǉ=�p�	�Z�n�X�:TɍAG���9**ܱ����b�=r�
m�S�:I��@c����ڥ���A|�e�a�N$����7�ms�����8����`�f���$��-FRJޚ���f������~4$yШOkO��e�ևx��b}� *(؀"c��XXQ�J�Q���?�Ņ��+�^��mt��0[CV������wt�X�g?�%�T�Ѥ�e� �y�ۏMk<�U��m]�������"�E����@�lr��'��x�8�p�z5 =�,�7�?L��f�(�l9X��rG�є��%,�G���' �.:�����_1�@ڳ6�����E��`�F�3LJY�Xe �ۜJY9���zEjd~��^��MSn�^P4�Y���ȸ>��#��3K<�*���y���G	�?�}N�z*26PG�ٻ��,���1���wdgu��3��E3G�{�L����uw�T�~.Pv�DM��QU��,h��S`q�c�t�ZGX��'��M�ӂ3�m65wH�$PZZͨ�_,�yb_j-��@4TFG%����x�h�!��]0��ؕ6��}�^r��~W9Z*�V�����q�/Ո���4+bP�����M����*%u4QDϸ��M�4p�oB��t��6�#W^$' �O������4{�%aY�̇7�u���K��^���ms�p���k�\��@�J.6��A^��_��Ϻ�ִ����5�=�
�3�{�NxuN�!�޼��Yj��Sj0	�#���� ���Y�l�en�pN�@�t�(�J����%��YM\�����Q`=$�י��@������|�I�dC!��( %RY\�K��)?�gd�2y®L��W�<���MJ4
����ĕ�T��Lh.Ţ��X[FrK&RE[�-\[nO�h��c%�إK�����'&|W�萅�F+k��"�e�J�2���5n�:�˔�\h|�]ڛEU�{4'Y��qE_*nvh!���I�g�̯݇�/�w/v{WFH��R�8��D�U�_��ϸ��d���,��&��{�5>;��J�������xG�*,�s��O�&1�>U��$���yT��W�����A��zC���*L���1�O�4(���#�f�S��Ў[Z�䕤�p&�\<�g
�?dZv*�$Ye�W7i"���Fɷ:,i�]Yl3��T"��rYͫ��'�pp�y���,|i�i�y�<V���3��ٞV�Oy���W8.k<����׸�Ʀ1CI]�&Eb-��e��N�+������C�,`��	��6#�xY�n>jG��(�^����+�S{n�nb�A�y����Q��9�e���+�APv�ߪ{�B��Z����e�l�P����=��B
w�:�!�X[�ۖ�:�#���@�:V1k���$��`?��\�0ə������+4Y�[�����0�Ÿ�m�KI�4���6Vj���Z<ͯ�Q��E �7DL7�?���44�Č�8l�%X�D�"���:�J�ѬǸ�a��l$!t�	�@=|G/>J��-Ĥ�Q_~��6�U��%b;����3 F~`�Ņk���̓�a��"qV)Ʋ��F)ڣ���
��<�UĐB�)5�l7qT�������g��O�2g�>+��O��z�(�[���4*�%��kt���*�d���~	@u���x�M�_�fI0>�d o���-�oa�e]Pd���cQ	̎���Q�9�����G�^�~켷_�j �.Y�-�[�����O�r�����&��j��{�����s���T��)-������#�Rf���*�;\�w�[uY]g����I�7R9���fཌྷ��#�x�S9�حޥc��$YΜ_�n-J���=:����<z�cYbf�G�B)��^.��� Y�_C;J����
g��||�� ���W%V�5��G���F�f4&��i����հt&'��H�2�ዥ._6%]1@�v��
��x�RPc��ןu�<�Fp���k!4���{Xl��ӯh�Ӝ7�n&v�uJ���!��qa=�BΊ0^����	D��v@�׊2|zq���ڜmq(� Щ�%�A��O3fYgb�Y0�*��-�/��t�[Q��(�1�4ટ/���,tu�џkhj��5s����ǥ���Q�������?�ˢ0������F2/1c��N���[$�j�9�Rs.�l�j��!K�B�S<j�l��1/1�z���>Y�~��?x�Ѕ�>��U��Wm����Ob��S�����n�4I��"ԔI�
� ���E�G��ڪk���Uh��T}K�[9�s[bA�t
MԮ�󏡂��A��Xd�G�Ny~!Q���Z�Z�ś�2�u��JQ`����!��xACi�ڰ-��?��TV����+a�M�ie��ui�p��k�M��0�f;퓍|=�- �HC%봊��a�w'�;���т�	iwb�c��I�[�۹����c�k�耵��VCx��:��x�gs�uV�=����/���sJ=
{a�a���Ie1�Ekc	.�ȣF���Z���ٓ�O7�X�-RR�����	�3M��{NI��!�m���7/p_Х��� G��\�i�0D�#�m�ټp�0�_}��a�;�i����e4C�T��7����J��e�qU���ۅ �l((%p^x�KΞ���,"1�a��Qu�Z�XbNm9���H�:]:j2�D>DO&]�@�-�莒I�J8�,���eL/�~�ͣ��1�ɻ@�o��r�O,���>�N_E��a�?��?]% S�0** ˪��ni��䅠��ԏ�79�c��L��Ϟ;�2s
�$�۬=V$��0ZCM����.�J\�8�%8�R{,��8+F�w��(?�7KNG�k3�qx��Cu�Qv��ڔ^M���0ʸ�U�H�J�u�� Q�U�A���N��ѓL%���f�k����b�K2Ū�Պ�:��o�	���mS��Lv�՞Q*�s��hjVkf��T�M��l��Y�f.�t��A��z��T��S�Б��`�����e#��S�w��R��O��%l��T��E���3[�pXO��0�P�X���9�(Ġ}X t9���*ǲ�\ [��9�8�T�V��ɒ�q��]�,��|$]��|j+�.j��l.n��s���֖~�R����"�"~����Qsm����
�Ӏ�(*DPx&+�����"�\���L&�s'T�@�ڕqje�����G�F��f}+2�56����n�I��Os��tC��4:���R�=7���B�F�{�$;���X�.]���-\�R�+>(�,���C��r�Q�D&����`��& ��� ��Wd½|��;>Y�ؿ���`��c^��חY	Er0t��G%K2��vt*��0F��9vɽ`W�Fy_��*⻼��� ٦����(f �싐��q2���)�7SA}q���'0^z��>��a��eaݾ����� _��.��;Lh�V?� m��o8(�Ia݇���v�"}R�B�57�S��e=�媆�ƴ$�,���	9�C>݁Q&�G�F�IzO��6�W`6
���:5iY��P]��ĭ.QD���y�f��_�>7g��2U�ɠ�ea�iN�!<���^��aC�Z<+\���[��U�B3���l��({S����DJ ��t�qV�	d�U&�k8<%��_.W�������O��r�n�KZ��T<r�c�����+]�"l��͖I�]w�o��vy�ީ(����׋P��Ż+�����1�7#G&_T2��
d�hJᢝ\�r�-
/����	5^��V󄤃q����=F��Wa#��!h���|��,r�=���]��ug���&3�!<�<�_nǷ����pTx�rfj-64�}�������Pʷ��obU�U_!'��Q���/D���ҳ��A�C�d�鬬�j�~e�����L�հWg�#�Jn���4��3�NJ����g�@r?9����$�,�Z^�rQ���QaY��宰�G�}���Q ?A%�p��D�LN�=���JC
E�ѕa3Hd��(`+��`{fA��)В�I�sIs��Q%�F��[-[ ����!�Q��$(E���v�n�"���Iq��ĮcM]�����;m�T�\q�X�L��F���P����b��_�ڃ@��S�k�+�x�=�ݕ�X��)9Jr�䦩y��-obp�۬�&t��l�kH���>���?O���~������7��S�����"�.OW+r#��Z��8�z�Zy����
�k�Sq,|N�C���p|ZD���Q����YJ�^n�i��	[�Ty�9�C�Y(fRsx3���d��������'ʎ���X�T�o�5����h�ص�(��оM*��!�WÜ���g[�A�cX���X^����Z(�6J�����S��M�*�{Y'T0��M���%�ו#
�s��6�cf�}��H�L�����������lS�\���I��Xg�X�� ����Dk�*�)"1��^��D�-�z��.k��@;P��:B�����cGX�h3ާ{ X�� ���i�� ��#�JĞ��E9�VJ�m���DN�^3�o!+�aD�48�C���%9����K����8�u���8*��T�>��I�K���Ό+C����#�o����>o�2�X{����}�Fu���W�!�?�x*P		��?W�6�\�xШr+�6��;;ڒ{cG�^�=L�{�C��G�7�8���Rw�(Cy{A�pO�>J��Co�ˎ_�9�- I�8Y��z��AU@�o���o���F�L$�R��	��wI�[A
�=�����5��h��C
�'��T�W��$/91˭�e]}�?h�e�oLr�rBt�U�H�0˘U��ّ�&ѿC,�VߝX1���]h��W�� �k�`���ف���|ܖ%s\��R,��iP�ld���=M$��"����^r������%T꘣Il��޻�pݺeG�FrN[���܇}����I�>�`F��@� L���y��	�ij�O+���Cv��\�`��[����#k,��K�����`���-��|�ڂ�1�#2Ⲽ�^��)d��)����"���ƬZ�xt{�֔y�B�*��V҇�����H�dmU� �1�%B�wI�~��Wΐ�Nn�A���/侏�'�v���6�j��W`�A C[�z��1�]��b��a+�7r�pϭfeC���ڎ�6_�XQ������_i��4��~'5�P�����A9�s7v��@��4���X�����|���-x���z�ԋʊ���Ħ�^�v�	�:n����W��*� ~����Кu� ����\�_Y�1���:�-��$���D�'}���u{�w��y�蕟à(�v�Dw觥�dn�`	�\�IڸG��p�������,T��u4��\t���:N�����pkG�H��Yl"M�H�$޻k2�e��J����ܐn��'���������8�\�M��w��������ŗX?T7Ag�]�%�@`���'���N���9���v"�m���U��J�/0���CH4�a��Vy������� ��I�}�ݭ��Š���JS�dԖfgm�r �>Q*�	��[�>^�8Iv�s�;۠�aA�_eͪ4�X�E&��Uv��W��{��yak�!G�!����Gݾ��v���O�
�c��"��_��@:Q����ù�Λ�x�K�����Yk(��;p��D^ɖ�m�r�gv��:�>^M��#���nrnd�]��ڬ�����Q��O�qw���N��R���?UP���>+��o�ڋ����OM��?�r�|���Dhy�L��1���A�^�.%|0�I�X�%B�&�eOǵ9��U�K���^QM�7�W��A��ܠn���"��CQ�}$�)q��o|� Dc���]���Ħ	��藵�o;�.e����GY�|v�J�� ���A?��	_�S���;A�h9�KL���aBl��_�W�]9-���ϊ=Ї�Nv��-�B�E�o˰�y��'�kԜ���u+��._�G��
�)�F��)K�W��'v[ƙ�6���z+5�q;�������
@�c�K�0�-5�v0h��'��O3JN_�N��/C.�D�St�}�<�ú8�SU��/������|�`�Л����l���k	�*���w�7���ؒ��95,�>:�W�f���-�;z$<i�0� �B��R����$�R
�!���ye��@=I�U�� �En��k�oN؉�T�K�_:�ӗ~��*@��b��7���0$i�	$���#6\4����/��"[++k�i� �Co����_�{Q3����m2�������bG-3�)�ԫ|�yoEL<?�7EjݺmAE~�� �5��v(V[\,m#�z�~e=L} ��ڎ�G��	�)k4Q�HK�P�t4��TK�[�>�t:��shS�UD#��:_�3����C���83P���J[C`;����τ���.�S<��H^*�N$r��z��-��ѵ�Y.�n^AaEΟ/T��M�_�h��4{��R��==
e>Or�$��b8,a0K��j4��X]�L���F�(���*Z�#`s�ɬ�6K)(��i����Ɏ���+R[e�ϊ��݆G�zJ��=t�-8�l��c��:2LR��tp�Y��p�mc�3ܖް0j���m!���P1�'Vs�Bl%O��0��!����A1ۚ�Z��ip5Wa�BG�����w����
����-�!��Ũ���Ɔ����L�Y�H�Թ�S�'�~eE[���C/$��T��<U\~��X�?��%��L6�l�e[�Z�B)8��ecuFIoq��\�Z�7���d,�9�`��l�Ʀ��Ddui�Ե�bX*b��?<y(��b-
U��Yr	���P�����/�5O"��7����_��3�0�G*����b�8{����CX(�B���dBK"��Q-y�@X�s��F]U�%b`���G}��V�"�'VP&��S�^�*HWNyXa�9����xܞ(���˩I��/∛X�/7�S@�b'J��M��I뙫7�Z�r+�0d����0����0�R�<����OAe���� ����w�@�t�.�����|�n�[��95�"S�np)�abs�Z��=GJ�QƜ�i�:�֫���\�/���1�r�^�P�Lb?2�*�h7ZM-�u-�|����!L�B�`�"����Z�z�H�$�R"*�7����16���(�P����.��"����hԀ�5F$��.��2���C��냶V��w����p~f�i�9S�8�U���܂%�
äG^�?���LK�uN���NM���V�NKa������n���u�i3M=�����@����N�����Dy�nR�t���nj�c�����Uc�9��dHa�F���w�:�}��4聯��`�]<�����9l�R�D�O4Ws� f}��ԙ�)���L�`��2�@[琐�O(p��E��)��5�U 01&�0p�lT��!I�@��8�-g@��!N���-�T���t�1!��!�e {�'�ȗ�ӫ�dr
񤞲��0'��d}�n�b�t	��ѿP�>)�A�	����eQ�{��xz>h�jb~������ʷi܁Y�nH������Br�7vN��)���{��W���#�[6o�m!~o#���}����U(U{��P	�-�}�G�T��j���l
V!6�nsy�a��Ps�,�iG/mK��rM�D��(�;1��qNv�L8$��s/�a+�b�ZT��ڵC����D��tڋ� `����!��� qzj'���Z=���S%��c��55�I�W]�|2ο2��$C:�W����R1�G}7��OZ��X�F̟��
���m���ѳ|s����Ֆ2i�k�K!E���ǣc��p���j�I�C��ur�����~t�]F�Ǜ��3m?�ea2	�8Lǃ��8�<���e����!��ǡ���O) k�L����$z��䨔׳]�h�T��|�$�!1�ٷ�*���X��xS�*�����[=c�N (ͥw�����1�ml��@�= �.2��5[F�*O6�.��������]w8�s {��I��	2^��o��� d3X!	jvN�2v�>�R{�S~�����1=O�?,&�k"��}5y�Z�@�?�4�1Jtܯ�S[�=����H�చ=tu�I�wzɄ��#���wn��  =��g1b~` =?��^� �>v{@�����e#\]�����7��;l��BP�;�5\'�ަ�F֌�C�����^�z1�hG&!�����ڭP�n�u��E����c�|��oV�i^i(�>��.8�݇�Z����iJ7z�&?x+y�{���8��n��P,􂥴�:��3\{-E�[$���:^B:2��Di����P��3�x��ƈ�%�?P7�gO��u���8$��]*�(��餵�0��wԑĝn}�� �3]-$�9$�],���&rw
�&<����Z؋��)�Jov$SE�3� KQ��
�-3�bx:�ي��_TG�$X(�%�)f�u�SI��������4͂�~�hm_�@���I�#�I�.#��(��w��,O�Kb���	��0 �6���� ����Np��	CH���	�~~
�@���&.��A}7��)9��ϸ��j�s
�X��D��4};�������W�{��5�p�W7Z�LO'�aρ���&Nf�L�Ɂ�?0�l��H(C� ���RC�m��G��mr,mɤ�V�0�
j5���cL \�~X1��^h �,G���Y���nN�O-�Ȁ���*��~���ݎ������W�`���\w)o9h���!�0ґt[0�:9����"�ð<�N����J@`ưΙU����<�_�џ��ӗB�E����k>��:v�~Ɂ�G�Q�����Ȳ��o��jvR0�,�ǂ������.}�܃|�c�`'7�zB��-�����S��|u��l��;H�AK/=ix3�#�A��7��ǀ��4��V!VAG:3&iv��h�=M=8�(��y\����Hi(�q'7F�0SG�i�;���U��K!��M� X��~&��"��.0�
n������|M�����b�<f�N��4U����7xi�X@� ����Q�Gr�"ȏ�;���X����7�9�U��o����B\����Ft<c�C�������9��%$��� �%����΂-��M�K�M��
![���>G
��[4�A��@&����oC��С�
���X�Z��c?,����s P	6�J�aӳ�������}@uשT�	yvf}�86�@�e�VR�'Mo ��$�y��S�a%G��/��UP�z��ŸS��u[�2�:�_x�9b���NCo \1�����p�)�x���R���r��������R,q-��N�_�9h��22@�m#r���CVU�²�����Bǜ���P�a�*r�2Z��</�^M�LU��֪&�x��"���f|��$J��D������k[�8������[�G`xix-����� ;�"��T("}׎��:�`�qg����dU*��˔E.=G�
4����O
�e�_�߹]����?�k!�k.	��m��.,g��e�emCz�8$c�D~�B���1t��!��6cG!�W�".�j/�q�ʄy6i[���F�����'����}f�'��אuǥ��#��A˗L�-:��!%��Ζ��M|�'�u�պ>��f�=��wRۇ�(s�[�q7����p�=?\�_8,��ĕ�۰B�l�PE�j�����U��aǁ���1��~L�B��ivx�*���E?��:��vA���I0�l�}$RA(�%_�5z>�$��	�W��W�ԇ��*��`wDGI�2�"O~���SBc�z}<اU�*&��Sa�ͮ=@��N��B��mb"�&'���F�a�}�'":,�p��!�7�u]M�Ü,À\�j�����֤Q�'��Ĭ_{�9�D2���/�U<��e�߃���I�:��"/4��O�9�U�'OK�����A�2b�tr�_�рRY.u���t�p6�����=��}��f|�mN�6L��P��Qa�u?#����Pe12h��\����L��Y3��K/�%�c\7I��y⒝�5O�5aR� �%9��=դ�JvhB�$�y��g6�-�`����,�q������ 3.$�z�P�q�k��G������FzAFe\��R^o�i,%������� C mQa�Y��5XEL'�7��@UDΘs2W��=>.�G���8��F��\1P���j��:U��Z���	�n��ڙ��=����돝'��3V�_u�i~�?������Z^-.˺��F���L�K�eAZ%s���`�,w��(k����s��3�x�n�v���_�8��M--���ΈQ��t%+�������Tu B�kX�t,EK�u����R�rW� M��fb�.+߷�Fb�V�KQ��s "�2��]�P3W���-�������HSu������V~��倜��>�~d>���G>�/2U��М�"��J�e�C��%&g�-{H�V��R֚�`�׳�$���ZP#*4�iM=�x�"x�r}X�� ��8W�qZ*��cي�dH�ih���Gl%���S+5��?�w�G��L�����|$�\j'��L�,�I�	B�~�y���/�9�&�>�Z����|�幏d�S��~?NH��9Ց<=2/��� �<��,	�>�o��Hu1��;=8<#A���U�:�Û������������!Q����
-u�1�(Nm�I�g���tN��2��7�$I��Y�R~l���LpĬ�~�Wv%Ok��u\���!Ova�ȵ�6���r�9�(��_t��\�ϭ��dA���꠫�)�H���l����E�Q�-l������M.�����"퀊�*dt�ְ9���>��4�y���i�Q��A�2!�$+d�~*+K7s�$�d�C�y=����A?�}:��ND߈b�����8�f��9n G��-��f󽵇i���a^��=���sW鉫1�ߴ:�K ���JB*��:q.��M7ɡȥ=�]�S���Vh UU���k%Ёx�@�P J�l���
�� �k�� ����d�҉�z8��Ã�
w؃����҃DKY��S�6P��>�}��\�R18:e�K}m�~pRX���	�"e� H��v"��>k5IH���'%�6N]uJoW[hsUD��C�dtG\\�����@��Mb{��9ב�Y����'^�am��d���N�1]�[OZ:޽�i�3ͳJHf�����B��ͮ�H��mA6h�����w��Vd)�E�;m�	J!�u�Q�-Liԣf�'�e�^�����5�i6?<����E�W����L�.홭�>�����М�&Z�ȍd������EF����"���$e#�Y+��풙���,F����:5X�~*/hYB�\�#	ո`�;~ C��ܫ�����8��U�p��e��K�	�H/���
�����u@[�X,����6�Kr 8#��gzǰ�ۜQ]��[�GٯE�9����c�"�wP�a���랍Z[�����)����@���}*�Q��w2�~���K�>�Bi4�uv��R_�G 7P8�����k՝�Xˑ'`�g>��YV�2T51�����ɏ��f^����g=m�J�蔟\����5q
{�jnR^�ڬb��<�P��3:������_cM�ٍ"��g+J�3G��I7��6�vI�e�!@�|*��e�Ft'H7����:��O-0ѣV�MP�:�:���?�,��
�`�[���_�_ȣ�u�� ͉q�ߩ(��T�0���ʸ|)���������y[zZJO
��&�rP+���x����WV>O�P�n�=V��^%�5Cg�~��� ��"��[��cu����dm�t��d1[PĪ�μ��M���Y�B��B&&
>oȁ~9�q�C����f������u�PE3��k�h	�7_k�n��46B�J�g~.�W�)�8vߦ?��[>����EK�mM���N�,�t;n�;W��ܾ+ke$���2:�W���I��c�婋߻ Д�+艫��^��qU"$�Q�>�Q�.��*�g�R	�}5Es4_\u�����x(�p&Bi����ڸ�������� �f�Wι�#�������x�K����H�Q��;�'u���F�}>'��N3��B��t�|䯹d�z��3�
�ћԗ��{�l�=�3�4�N���3��0{�|#��M�e�U!�4�B���?_n�a�*N}����.:Q3�疟�����9b�P���Xm*���� ���w��tib���~�Nm�d�V���#Q���<v
����Vj\�8�SY�*>3�+a����\�v[L��zn8t³�\�"�+��:�&)B[�l��+�Ժjl����y�caL���}E`��k$}D6_ڧv�65:R��J~� �$$������Xu7,�?O�oc�Q�Xd�l��|;{o�i��5&2@�Ɖ;��>������[�������a���]�k�a��(���A8W��JJX�R��[���ɧ=�Z�
�>���`�JL<�����ɜ�S�Ү��U }�1m94��<ܷK����/%����yLJ�k�8����(Uޫ�)�p[��e@�������B�/v%FE��0SNM���;� $�v V#G-�^^HQ����Z�X��*������8������')A��L-�d� l! O|���l��Q�#�UMgK����,��\q���fo:˺a0S�	�(~�a�{�*I� ꉞ�ڄ�ٰ$8��RZ����+>�*^y�Y�Ѻ�r�O0d23)9bo�ĥ1��1>ĥ�l���َ,�������e�g_L