��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��ga���<�\��J�ιϛ��%����EuI|hV��H$�y�olgl�r�5��a�y�ͼ������N���~�8��/Z��!K,��=�Zma��Ͻ�>����V��[�	�|��n�Xq[չŚ_�2͒���2#�=8��U�2y��VV�~��Ì�a��h�5�;��3u5���A7d�� �Ǜ��VLuFM)���ө'xU���ه�Fk័tR���[����B5���C�ˊ��f�!����=�O�G����g\���v�:��T�:]��ξ�����+���Wc0�x)�+���yt���ʘ�hYp]����Y��h����H[�~yS��~�S��pX���O�8�h�km|Q�	둶}�<�������Y�`}σ�����t.<�|��;�;� ��B�A��a�����,?����y��
x�#`M6xGA��,$�st�8E�G<T��m� i�0/P^��msh&1,ݎN:�pAvf�q��F=�]jmMg]j2���%�&�{��2-�4m]�F�Ԇ�=����V�XX�t��ȋp�lȃ3^p�1c��#��ҍP��tL�d�Wd>�Q����aqݢ:ԥ���E� ��X�v��&@�h�᭿�0E��P���]\h���gT�9�Ɓ0���.��P�� ��p�I�W7�|��NAr*��>\T�����߿ ��Ȫ����� ^�
�K�-ux%#`��\�����[=f��G6٣hג���Gmb�P(����x�@�NfA�\Bհ�Fr���c�BD�X�^51{��<Ҧ�)�Қ�`��)��-� ��6v�J���A:�K0������hA�]1 ���:Bt� ��������t`�.?�ƈv�( �Y���*�q�L������&$�j�O�7M(_��-�ˆ�B�ꉹPMdR��u�
�t���2b08zw��2l��h�μ��~�N�����-��\��m�������`cuzNT��Im,pʅ�Q��|�,p��ߔ�K��l-�;q�0��A�~�H	�r�MNj��w�[�z��QC����B�;�A���� @=)����t~�Q�U�?��?��@����F؊� Xq�0�g��,�~ M*�|���f����-W���rbw���U�=��5�o�xk��`_�C�翼h��Ć���������UN�E�[��+X�[�5=m�s�)�:�+*�Ux�����}�S�e�ƈf��#SM ̋�P�8�BJxQT�e��;�I�T�!�r�\�}P�fY�k��k�����?R��3���$YfÅ?X\}o	c
rHE��J�0%d����C�!}`H��_��"�O+XOʳ�\�-������o�4�̻3�v�%x'���%~$�Z�d����âY����#i�|s]�����CW���2�M�s5�dS`1fB���N���I����'�tw��/`��J(�>%R�ݚ��P_у�W,�^z�:��5��L�arA<����4t�����*т�ᖭ!�ϧ�����C@�\�=�N~��hD�S�Sk�P2����Qt"��~����S�����KZ}��ڊ�.���N�ywl'W��<��@3X#������s��
�N�����������ߤ]ʋ�%�1��eqɦ-#0�x�u�`h��
6r���_"��I�'��Lx����kW�g_dq��G!�Y�U�.�>�XM9�V;WX����\Ѽ&�kCA{c(��x�����r��xg�U3����J�Pq&N�ccp/�	�LOЅ��:�\��J?#ɪ�uS.�q=!�9>�;م�Ӯ�F�qE���F�7�eA#��n�
3��0[b0��
�������'�6.�a���������8dΜҮ޵�I��;CPRf ��Qa���=I���е�K]��n^i�٥*v�=��,oiO2������WZ�@��&趠�%6jr"�2orhAFR���-%<�,��J��G��Z�d���R�D=%*��p#��!���'�𖿑�E�Г��;��N9~e��xen٤ee����-7����u�XȨ�b�wia���BAI+��i�Xh���FG����1$�\i�*&�'� ?�!:{qQ=c��7V8��e!�����!�]�_���k���s�QK$�m3�_ׯ�hn�m땮'W6,<.�!�Tt�է��.D`������o��GRi��xm�:!�g�d�(�\0���&)~Ӛ�UI����E4nb�����$�U��A�v�T%��E���G�Z*�<
?��AT5���ra�duP^8�� h��?V�+	�]������Nծ����Z��-�����?��<�6�M�-J��k�'<`�{l=I�.=�5Q]U�-����G�`E�%��q��Zs���MF�O�9�~Cn4c�9��{j���u��h���"M7�yzǷ�F�ڟ�БvF����4|+P	�Xu�P/�Qm�����;���O�B�m!��)����A;~2q}7�a��?lU��	�c4�\�4�{�?���/!����K���"0�f띃���:mp0)��9�:�>\f� �UU�����:P#���~�e�*���K�d��FYx���Gu [քb�b�}�yĭ��|<�e����C��w��4v���S��}�3)j��'pD������70R��[pE�R���@>��b��.w�K�������xT^����WlI�-wi5��%�*'���Qp�`]�.���sN�?l������ )�:��$������m��;6
^�n�Y��$�
���!w�����o��h<[�8�Ll!z$�59GA��-Ό��[��	ljC�x�p��G�8Dߟ���)'V���D�-�*��b -K��[�y����5 �K�u��2J���@-���f^ԚI���"�E.���d�&1`�@����ץ�oF	w����ҡ���5.Y&�Y�0.�����D�'<Yz�M��է+���xL+�(R���غB`1����J��ݛ|�ÑOqW=�C`8�A���fAw%=�w��B�[ <YՔd5D��龨׿�������	����;uU̝��� �T�@�$j'9ex B̛���g/s�!�M�I��o�0ˋ磭.�T���5�4	Ԇc&��GE.l:5yn�"0i�J'8Æ��A����?5��5�V�:�Ǡu����bÔpF�D�6����=YȎ�*��� ������%��E����V�����eJ*Ï���a�i�/�<�'|"�������z����xy~���:m�}|�*f���(��F�	'�|�}��%?�S! ��+�����9`N�p-+�7��K��Y�z_�6�Z�E�{JY��,��*R����F���V@�5��y[�m����(���|�J���ԋp_|�9E66���ٗ��m�^�t���3�ȹЎsL�^��fyg��	7nT��Ӧ�|7�O�����,t��|8`H�\JP��*���n"/��P���� K[s C���5��s"ap�ƇL�Oz���zC�����1��X���؊�A��k^�16R�y�5�'��@]����PX䮆5�,�F)����Y�ɸ�[� 尵�W��Z�c�����!G�$h�5�x8�bJ#�2"���o�]��H��VT
�G���ҷ�����
\#C�B�����%��S8@���wL| A�|�^�#D�3�䙢M�ESo�?n�T����[���/r���K����cvnF;��|S�l�F̀�����V#X��߀Bb|�Q͑�Gi�b#��X�N�F�J����j%�GC��%3r��)6��eߴ7�����Ç����aJ���6A���r�.�|�M2@
E�������&{�ǽoF.&�����*�v���wV��?�kՕ$����aU�vp{3�9S��-L�����Rn���腶CË�;�&�����.�� �!�'s�Kq�r��ĎM����5����|�.�����KPS��E��$i�"��N�hCt6w��V�лS�q���{2����˴�=�%K��:S��-�Xq�ʧ�9����iO�1' �q�l��96އiy�z�O�����7e���E%�t����Q���[ݛ����MK�$��e��u�&��b ʞ�-���è�&>�֧�y����f�2R���`��	B��*�<{+�����n�]s�#&~���+�\�������Q�4�����'��7b����1p�%(T^�����_��kZ��R�iV,������kYd�	�ۡ�.�_�������P���l�kа���q��ƈ�3���� wɦ��Yw��L��{�M�&�B��<���}����`+j��W�s��G<t�"�<f�Tq2ƍ�2�L�J����%�z@���E{
�V��RŘ�ûЇ3#Q�V>��ڮ���k?bɿ��� �<Gc��>��L�����Ҧ�y�P���a$\@ٱ�:���d�tr�W੶�GT��)�}���_�촉���4��aF�o'�H�Uy���m[>��7
%:Xc��	�~�Ka�ϯ���	d��z	�|8����׻J�vv��D04�5�������?���T�pC�D����n3>��"��=������ǣHؖ�t�Ŷr���G�Ye!���w�E>:��������ۣPYZ;w޵+�N;���`�OG_�Vl��v���#����߀s����D�Yf �=T��\���dj��X{S���S���&j����W|v?�8���t����j2ơ�E�\3!�n���@0���;+�x��j�dT:�cN����F�t����~b�t��LO�Xg��/l����l|��b`ocHF���1-r=$YD]��8���rs9;���:"F}e�ۆ����������k����*6��ܧ�6_�,,�pB�rM�z��r���/ǟ�g��Yl��M�˳w^�m?O�*��/\��KZ|>�9@A"���<I�����}:oA�E�#E���Xy��R��l޼�lD@t}%�1�'lcn��b��d���<kX*����]��k�����6��r GY����W��
~ي^��V�~N�Z[���4�$�k�&���I�,S$��8X�ڠ��	m�=Y��c?^�����B0��}���;����Hw����%<ꄓ���m���]��~R2��� �3<�8@f~��7�XvW�6�/�*�K�za��e4#�Mju����94�Y`=�#��&}���=�I�?ѫx6~����T�q�-�KBأ�O��ǫ�X������a�b���^K`'K����@10���@�}��}�f>jp��_]2�8�?�-��'߁!��T�-�G'~f|莩@�U�NEw����魤dT����ϑ:�v��Nj�ũs'ts�����2�H�WW��w��e��cI
r'�QPq�	0\�5V��s�Sm�X�ٽ�����49�O��Y�k�#S��vjv�7!vV��� C	p�m��Y�4�C+*�D����{�X	Nf�Ļ~�G��*L��2P��a;?�L]KH�2/��r�΀�C�0w6���l �a�4x�q�w  �<�[�����m<����2v�T@��G#%���^6Tvɤ�5��=��T��[4ۯ�P��J�ƭE��+�6T����d�*kk�p&�|0���#��Ctwv�i"�b�3-C�St{�.�&��F�eE����TwqfU�4	D��g௮�g#�b:�z����x��f�ʉM�������Y����|��S��&[�f�JA��Ä�h"B���f� �s��4F^JӴ�a4�fE#�ֻmN1g2�T/�H�X�\���,$N=�O�s��3�TYV.eEc\���A X����0�Y7� ���L~�oN�� Ǘf��JH�"H�U�#`yw�_w/H]�X���2���=._���{�;��c��N�����&Q��if��Q�:��w\�Ka��lj0Q��q�*0��%^��bO�?���{��W��RJW�u���E�蛝8��o~�����ý�5<6��
� ��s_c!J�ܹIw/�[Y�r�a���O��e�n�ʮ�^�Ntx�i9��W��ʮ�а����d�k��F��ܘm�䒘��Ǵ��E!p�����p�4�s�?^
����%�y~
�%��t�(�f8<��S����)����!QWb���!�-ݰ'�4�>iY,�Y��+i@8��<��^� ��fw�8� �M5fW�^���Ҷ�t"��^�im� V̠�0tOt�y�
U���pO��8s��z�RF�F"c�w�H���o��
 �Ǽk��%�A�l���#��|�����9rE�N\\�����E�_@�=��f\��h�gPvJf"I�`���jP� ��@�4��Z/#J�����ԝ3̫�VH%��*-:u=	�W��6J�U�[�^KL=+R$������ݮ5à�ԁJ�g�:�{B���i_�0��z��K�h4Z�Z�o�
�a���7�C|���{��b0	�E\b}�ΑF�rZb6͇8!P"o%
���͊I��)Q�8�G�r�Ʀ+��F��J���!�1/�11������w������ì����I��¦_��?���N���3Y,ɘ��v��ށ��J�c�0��$=��q��M7F�H�����=h�e����O�/���+exa}��$�95!��e�/:߶�t��jHZ�<�e.ҺHr�i)�b�����։�'Q���d�\�{ q=��-;h谝�5���\=l��yfi������MXF	wC�Kp�O:<�$�C�%�5p�uQ5�3������.8��in�^E�R5p�_$�e�{�����Zll��~�>$a���g���x�k WʐƗ�`��eI��x7:�m^�	�<�ϣ�;�~M�/W m���@g��x�t_b�p�Gr!�vIȗ^���$��S�/A�:�-�a�I�EN�j���T6��8f[�O��+U�`�8�������$kVV�k��(�y���O��±�v3�l߇j\!��z�fz �xn�Z�Ȥ���5If����� ��	��9�T��8<_�#�F_Hwn�+T�$��_YD=hٌu���T�8��[K��V�[��I�*o��ɆX�3�@�B$〽9Utm���+'�A���4s��/.��ä/>�lX���^^Ӧ�'����a�t�mA|�U���"���e���l�_�����S�x�] ��걔b8{k:�T���ϲ�%�H��Kj1ø����jd��
��5L����H"X�6�8*|�/������M��+ds����ׁErEc���lȯ٧
��ʒ���KV��ўw�PO�f��I���0g� �;�F߼�
��Es�=T@Ƴ��=�Mv{��ٲi��d�	�Y���jD���Um��ǅ�AJ7�-QP��,��3�u2;5��|0�6�1Ou����Vk���4G��*�,���lj����'j���5�#n5���Ӭ��q����&ե��Bv�61�����g&4wϧ�Ɵ�s�	���Q+7��M�pm��=8٥�^�M�%Un�gݻ��*���D	�P��ɮ��  ��}��ځkz��@]�y�a^η�2�a}P��p��qoN��
�k�WJ=D8t������=�ɿ�r_�ۍ�R�E�ro��W����?��^�T~q�Zz�S9���2-� ��a1�l�t�&����گ���"ۧsó��y����wGj�8�YR���dO�E�v ���T
q#S�p� ���Z��^��U�3�����ģ��E82�^(�m����륎�{�9�$�*�܅��V���=�K�n�e�w���`{��5y�W��3B������ׇ2�Va�����_�@[��	���,�e[�P���d�������7U�/�#m�?�o�9��1���tܶUߪc>7���,���fT�����X�^������i�$���X[fܞI>���9&?\ۻBO��֝3�|c�,�����+!����l�XV��K~+tH�X��P{���dI��{T$������乚�Ś�l��AK�I�Z@�䤒:�4OǓ�SD��� ���(y��Au��eydбÇ�!�����ޕ-}�#�-���	P|1�!NT�p�l�H��X��~x���3$�#����x�,Z��!�sɣJ��D���9 ��js?�yP�3%g�z���d�ީ�s?5��͗O������B;r����#�\��A���B����O/��^�|�6���ve[x��L�Z��n�0ǋ�4y� �bS�J�[�m���EL�CB�_�i:��^t�t�X_	��C#S]bT�B16�<��dQ��E4W��-�����1��Ag	���;,R�`XCN�I�L��άVK� k�/5ҔRt6�v�3L�R��ӥ�Kˣ�^Ǫ>u�+Vm[�LS�W�} =]�B��
o�i�����2���+��Vͩ���\bP�V@��o|�ӧm����w[�,H���(3`��U:�oN�9�B�5FCp�z7 ̅�ue��r؋O��y=��L[��E�C����H~�8J���u��ǻ[߀��2�ɮ��%�f8.*1���'����u迟	�2�Vi6F�F�>�ұ"��/�c�k ���2�,BDGE����.~P�&R��u0�w�M�x9֤2�\�Ӈ�|}�rNN�oh�#��-
��U4�<FYU���଺�&h�Ia�����x��P���fCx�I�G%��a��n��}͑�n	�F�\�)_�xx�԰�T"�C��t�&�������������aR����.{<7�o=4�'#|��1�.�grhM����;bB�����A�y�uc6��E�/kA�^қ���ڈ�2K��z�=���ֳ���Sc5��y��V��.��6���	pwoW���/���Ĥ�4�'�ި8y֒�o�J���1쵗>;"u'Y�����9�1�P'�qN����L�.mx�}M�s.ｨ��h$��v-�_�I3 [��Au��3��>�ӝ��	��>lZ�	�Me`�ݭ�{�uU ���#��L�,�y�N�TL�?.,o쵺l���������;f��k��z�*����������0�#��η�a�In�La��.A[s��kcpgH{��F�|^�6���Ċ���A' ��O��bM����.���ao����Q	Mi,��5p�������Qb}Ӵ#Q���ٷ���/^+i8��k��|j���IGF+΅���N�y>?kH�wl���W�� 2![��"JZ���h�b�7���������yt/�K4>�1/j:Δ�[�gh��N��y�o��Ho��5UóF�x��t�����j�&��5��dI#�]����֖���0a�+!yyA&��B*��G���xw��l:����U ��}K
��>�u>�ٰX�ꪋ
�R����i�����x�K����p ��������RF�/,����s@z����i_��+wV!SUQ����ސ)7������{���c.ў�&EW\Lw�D-2�������
��aG�"UY�v��Eg��_T~�qI���>�٭�T�ӕ����=:���;E��	a������"��2���a�m���7՞�KI�{|�� Т���,�;#�g�d����b�5X�9�f0�,��cDÓ}�N'G邖#+���'� ��I]:�6RR��,�Ǜ��Kf� 	����aC���o��煃`��5��Eַ�ۘL,����PR��;>�Y��+�Gm�\H�!l'��
���;�S�N-�Y���7�T�)�(0�3&'�j��V��	�NHxVm
�$�x��n�
�����sA%�@{�?�{Y��a�*�����`W1����|���[V}��⑻}����Y�=���-��\0n1�2tl�/�X ����Sx�L���$J���hW�T�PX�����XL'�^=���ᩊ���'����Iٯ�$���l�}�4�o`���2��y��n"o>��ywGa��|�ܣ�۲�5����]��o�	��NU~$`�r�����	��Qp�����;*�Oov�kc�v��&�)y��\xɈ5d���- %j]���ЪQ�P= �#�'���~��>� �E��Ht�F����ù�^����,�7��]=�� U�a�?�MgEFp��xt��-Ran7������R1��RKc�ar�,������E8D��Aْ�&��m�}�bA=2�����Wf0Qx��������|*A��%�`̸�A+|0�"'���k������g��?�z���O��}%F!X�]����[�sB|k�d���B�e���������`@�O�v��ʘ��2��t�^!��Z����\ ��uS\Cl=j����x��f�K��&?���{ ��\�9��sP���γ�.9rb#o�T�'k�=5@�!3pv���(r�^!s�=�D��l�=n�JL4&�Є���F<ϧ5fHܠz�GKKZ<��I&��>�F���<��~}����&ծ���� �C�!3k��箕�\�Q��%d���h�m�?}Ĥ��(L̰���t��4�$e�������rq^m����?�+ �ӉM�e��{��؆?��vr� ��q��S����z�:��s��o�@����I�S� �@�9��Ǿ�Oj��~�\g{5�1>�5
p!�&m Px�o*N��W�شk�t����r{�~�����(߼%�I㍓�Ӊa�Gf������|ؿ�9�e���0}�mfX������7���	��^I���R��S����l��4�LU�T���@�[+��<�N�Ǧ��W��Y�F�J�?�=�:�����cF0�{>���:nJ�$��( À�:�?5��	��� Cs�4���!�X8�)|���hT[����Ji�	�$��`M׺�:���giq��~�z)]���8 ���΀%c�t��b_���yZ/.̆���Ę���!�l�Ϲ�D��P�D��H��q�<�J×�0���ƺ ,�%��C(��j�W)��0<��NL,ƶ��$�'��H�v��C��ģ�
W�<���.��y��`��!�� R,>0R 'ۊ�r	_j����u��~�z�@���>�7[0$-u��3@F$%�[Y���A4 ��p��:m*:�>7�S���ѕ��3d�c�_�ç�d��k7%��3|�
)���Y�u�Х��%��^m�A+�|_{hC��N�޲#�'W��._{D��}���X>���}�k�^ҷ�<�IJ�7�m�%g�L�Xd:-�X얧�A�9&k*������h�/�.W�N�r T.�J����,���a_SU�a��`%�#M��4��\*1~"��C�GQ�/�`�{�QQ��eb������ǚ�j��������]h(w->,-\�LϵM�6���տ�y1�1�|�f�u��u�|�gP0 ��m�1�E[�S����(!)�A�d�zGǼ�yCS�vm�+2^	45�'A�Н5ƅ�a�V��H��2:��F��*��O�K�o�!vyH���r�"���г�>��e鼧M�>�������Z0�:U�N�*������E�f:.�\g=��J�%IeL>�;��h\�8,U�����EE5D�n	:�QgU������)J�РB���q�/����X�F�6{؃n}��ଋoy���� ;jz�&I� o[u���}7�%��d9�+�Y���BYhf[�^�H��,z�a}�k�	yL���Q� ��=�?���R��;��*0�<%�EW��3���{"4W{9� ^*��z�)G�`�*8����F�Y۪ᣙWJ`�M����xV�C��z�Vzn�5'S��t���G��u��6��
 R]z�������i���:�xQ)d����04��>��v�����Z5���!x!ÄxЮ�8Y�@B)+?`�zV�i�_�才���gKpdStt%,��)kM��d�<��!�lŘ�]�i8kִ��9�xc��s�i �����șHvSC`�:��l|�*Z6 �,�"�f.��6��D����@L��
E� �Q���=��~#��	=l<=Ή <4��KOu�a���E�'{؀�U'�M@��o]�Xzn#�a*oK�q�f�b/�b9�
�@س�t�j���'� ��!Q[p���t�w�0f@��"vZ���u����&���-R\��D��#����MEp��{�f~�nJ)6��PF&h����:(�&ş#G݋�G���]b���grK\U�rmo\�J�Y<��14A}Wk�E4�5�ug)HL��X&�}5���2��t�]#b��˷5�y�?:�]zѢ8o-,����s�EV���1w��"�����Ն���[t��Wv}���z�CQ'�H3M`Q"���P���]`�H�2ë'�մ#eam0�u���~`,�p�0k0?P��]�F�emh!g`�qYD'���}x�o5Z���K��x��Tgs�G���"����������,���z4�5��z��i�� �Ѕ{\'%��Ɵ|߮��i�����03Rb��L@�!	�CU�!�b����/�����*MT&��w��3!�	��e)��o�ǈlf|�r�a��s����)�i�(r��o�V�`�2if�a�q|vr����Ea9Pf��!�:t��
e:9OE���Pt�Q�0���*��!�wv�t���X�kO*#�x'rb�C�V��&�	���hV��-%�GsA���)p����)�1�?�ٗ�ԕtz��nV_q��ѕ܍������<����g���#өW�4�NVW}�k��=VA^��o��0��R� �`4��.��׍9��D�0��e-�b!�<�$��7�9��9������쓪���VxJ�#ZK����d��d����ƪJW(���m1�lHb]���y�aݑ��f�ӻ���#�h�\��|5nJ�9���n��e���b1��d;�!N4B�` �}wAæ�i�I�;w�wxu)%��lαY�%n$�'����	I��zo54RӨ~�͟4D��Áf Rx	���p��R�xΌ�C�d�3C�mL���6C���'ӡ��������Ϡ�A�ؽͪ&�u�8�\
OI�="��l�!��̟]u5�J8;9����!&�
t��՚bBKv��<�K����<��QC��^L?��h	-�B���z�}��>{*�`$=g���k���cx���?��YU��CF����k���f
��LyԸ��{�O6D���+����,0'�qx%q��_�w�KT�9e-��D�� o�]�:�" 3F�.�n���O޸"9C+��N�+�+����{6��:��Kmd\8��l�i�:J�>|P�Zv������0�*pʾ����)���_9ˋ}��+m���SC�C�_�5��_	�y�o_!!~��(�\���1�(퇏N\2�ztu�=�7��l/k��(.��X�����k�'��|�?<�Q�+3�=�3H1�a�*;�)����!ћ�N<��TyɃ[�)��+J9�o�!��Az�����Wt���+��X8�o+��g�t+��j�������N�h4m�V���`�+� ��޼�	���f4$�� Չ)c���܄f���ݡwQ�q
�I���3M<�ǌ��XB��a6,ڣ@��<��Zֹӯ[�P��A5Qb	���%`�f2�/@�]���>���2���虍�SJ"���Μ��)�%��&O�����v�v˥�d��~�L�����������6e���rr�	M�<�JMd�Xt��Ġ�|������� p��̤��mkX��n��d6��/��)&M�˺:,��G��5��gU�͜�=2td�zf� <s �C����,#%G��o6���υ��	 n������B0���3�P@� (��12�({d2l����4ϩ@՛��]M�`��|�^w��n��q.��KH�����e�?( �L�O�E�G����}�p3M��hL�j�
8��%s�-�׍mAnQ��@��er�5��x��w�#
s�.<�z��#.�2RW<����o#�OD�� F��)��&h��@!4��^�5��P��[��{!<8��]D8����ғv����=��%2}.F�	���-���5�h[b&{�:ɅWF�?�����wb)tέ��̅@�*�Q>+�# �p,G�Q]�A���J%�1
�c6�Mž夅�ĔI���:S^�Z�T�k�EM3ZA}��"�f�M��.Պ��g���]t3�^ô���W#HHg/����ka�[S�Bf�l
�w�k?��5�e+�~�^�Q��h�����W�@�eKUo]����]�Ī���>iǪ�"���P$���&4ΐ#�	c���r�+������r3���p�a�3���=e/�Z�69�ɇ�O�N�J�]@<)%��H������ �%,:O���u�-?;yY�z��>�y�����f�\ӕN��s^�J�2x����	rſ�	X�`Y�XJ�ǇN؄-6^�g�ʗQ�li�7"�&3�\R� &�D"�ڂ�o�k���094�eh��S!8�j�(Z�IISN�G�98j)��X���.1n}5�/FB�JTw����^u
��_h|�{��E�m"�P���ۗ�;��t�	��d-	�O�c�4E���A���]���H`���Hd��%v�:M�A�ˁ>�
�� �[̍^�4
zR���/Cl*���6�A����j��ew哽�.T��Y�g�csYV�Cc<\<Bi�V'P�6^�#tJ���_��f3H�v��i�s��B!�o��R�D���g����	C���F䪃|�u@�S�D�kd�(��팲PGD�y�)����i�U�M��\r�;1R��Tx�*v� ��Q��iJVz�t�"cyY��A�}�U]��k�ę1 ʊ`ܧHӶc`�Ro��ڻ��6����=pe.&��'��9���b51��-Wy�_c	��N���Eى�kU�w��dA�?�S��BH��~S�o톻�R2jbqъ�[D��d�t����d@��I8����c�ݓ��:�*����Pѵ~d��S��W����>�;d���������M"�(�&��}ڭ������_d+~��Ͼ�'\դm>�&juVhv� �Sd��Vn:���Y�"�a��`c  +h� �&��*��؎�||�kK6ሺYk�m�Վ4�4�}�����O���`�y��jw�9E�b�_�q�Ջ�,��C]ې6� �o��W{��[R=���.��A������9�p�O�vd_�OOt*�(C��qԝ��ƢV,�l&�����m3W`8��cO�A�X�FH��$A�͸�J"��WL�w�e�	����������zp��UT�_���a]E�Pj��>�9�N�{Ïl0�"s��A	��(�0�V�v���})}�3���,�0��[�/����5��� g-h�%"�*O�+yU*H_��o�U�e5 ��WZZ�@ȁ��=��hߓ�b �`�a��D��� x�D�`n��d� 
p�<�M8	�j9�QK�}��EN O��1��i>k�8'���W�HH��|�H�J�(7o��(��-%A�ȋp;p�����.EĮ��̉�����K��:������o�Fe}�ڲ������\����am~�D{�C6d�v/�تa�����>g�R�_T)�dRïL݄��Z�M׮ӽz��+o�.@�fi��L�"Y��I�E�,2I�IA�!ª.ȥ�M]�ˊO����w�.�]�ND�����<v�"u��k�"��}�k�!��Fe�,�lc�;)��n�B|IRY9 �N'}?�������RZ#��Q<�z"ٜ&�8jE"��m�e�كd*�	��IO�)
@=@e�&������� j�l�+D��_�S�#P/ҏ��L�ܷ}*���3<���Ǳ�WAأ��K�\��'u�L�;�3?��&k�ײ�����+��U�̺"8��/F��r��>����JK6� #�uZг����f���������|����2L�y��{��yN�C�d�)&�F��D��5ӓ� ;E�E��<<�эOtr���"A�=jb�\^+a$������*���6VV��5:�W{pY��(Q�\eණ���Ǐ�P@�{�[�D`��xTw� �~9Oi߫�*�>�-#5i!���{h���UiY����[EJ��z�]�ia��ב ��^�{2@���y�(&���T�����ᮜ2T���P�f	�/Tfͩ��M�GR���#�+Y�ʢ���e��<���S���M�錗H��(zujٔ�l�nu8���UX&�\��0l@�-/AT>Py�����8��H�o᲎��j���d��8%���{z�)�]B$;��{Y�������=1���,wE8~��4IE�5@i��, w����MD6��~�`D$�sـ�5�wR�H�C$��,u�4�y>�&�K�H6Y��A㿣%�d�J�:A�(S�+?�hA�R'��,>�X'�� �gM��h�+S-k�בI_��\�����������������Hj���gm�-�_ܖ��Tb7Q
UV�ݰ���x�=q.���vP�8�+�BV�D�:r��Um��,0�Xm9"�9x��[ѻA�����m9��%�v��M����%l'9��Xq�9�ɷ�j4�	m?����_�|]pg�\�z����zc<8����\2x��`3�1���y���i������$���?[�&����Re�8е�����/*�.�^��/���q�WY��Rܨ�N��Ǖ�q]��k���J �B��P�D"��w����4�d#�����#�+�f>����^Sob7�%�~[�)Br� N��n�>#���B���'Б�C�3y�史���]�9�l�X�6��Y4�f��<���!Mz΄�?۞z����c�5)�'��)�n�����bn�<���;`�I�BG�����gp��#Ԛ�{7Dg3�5!��*�>�Ɨ�]��<��\�F�޿�7���gS�3k��B�hX� Y(�cÁ@�=��/�������R����J���-d�;ķ"�p�3��o���1�d������nd���Ø4=vy��RS&���D�s�C�V�cκ��y�[z�/q���}tb��!L~�X�7T�I�ك����
���&X�$��A"�f��=���Õ�Wko��$��vޙ,V@
���C=֔�/5x-���w���+[ጊp�9P�3��n!��dK�S��M!�!d.��HO�ٹ�D��܁RAF�gg%�t"���|�u������r$K��F`
B�.��۪w�{W6񂫵�ڴ��O$�a\���aAl���e��u� ���W�s!C	�>@�%�����
����b�jL�ϫ��.�7`��(���Ŋ#1|T���� k�nĐ�63��<t
ɖ�#G�gσ64�	M�<��j �wº{�1�P�]#qk!���ˣQ[����W�����_��2M�%2'徰�^�~�_����Ȕ6v��� B�A�L��X8C7�������V�q�a�}]й@�pM~���Ӗ�պ�>
4�W����O%���{�7���[�Ռ���w/�93��R�'a���J�oH��G�����ԭ!f�ѬK[f�U�A͈W,��������I��	-�S��95����ȍM�v��?b�=s�s���PrypJ�����Y�f�/��4R(xMV�n������Qw՘Ts��8tIG+S��"y0�������&�j��G��}�PIc�<t�}�\��?"GT#�ʛL�E��+h���h���jꞢi9��V�D*8����¶p%G.����U��ZD���v�����FָBv��c��m�?@�&	铻���Q�6�n��ܴ��y��1{Uk�L'���e �3_鋖o���d�z����FSn|~��D7�����z�r;�Y�5�A23�5ĸ�ɥ�N�ਗvk���.;Ѱ ��<���w��i�r�E'DI��`s5��v����X���u�Mʇ&e���c���ES[ݸ�<<������E�gk��D]�{�->R�����V7��Yk���[�I�&)F0���*=�<8R�ʽ���7Iz�}��́}E�U���9T�%Z2�f���:�}��ן�^R�v�[�W���hv�}/�]a"��@�X�{�l0�E�lQ:��@��o��S�G�n�a8�@���O�4���^�Y�ws��~:�d5bZ�&O����.#�\����m��7���=+�'}XE�x�Г6Zg�s���1|@��f7�i��*[3�_��F�WK�u�Ed�th�`���mȣ5lf������)����L�A4��H�S+��/�L�`/��a,�*_�}�K�%�����1��f�&�m~U�C'��?w�-�(ߞh�g%���K�o�)�6��
y����rwbs(�>8��Z�w_h�%b-�$v���^i9Ew0Nz��M�w�eꡩ)g�:�V��izx�Q�����fH:�ǿ�a��������������P�;cO�	��=
���B����d�d"�v%�7>lìFܶh�����O� n�bQڦ޷'C���4�Ė�CzR���1;g%0�8��X�"��<ė��