��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��R�%��«��7�:���c#�h7�u��k�u?��V/��5w��_ziCa��l��PQ'O�	C���J�#nW3����G��A?�k�gĒ��t��r5�,F�ʗ��gZ?�z�Z6isG���ֲ�nm�޺�����)�C@��E�?���x���U�$��������	2.�O��˼L�踂�>
9�Q
�T�&��q�_�Dê��c���"��xN�)p�&�:�x�걾���[����"�F� ���AH�f:�.'����%hL-CZ^��J�SK1W?�������th0�-��T��K�~D��'�2�9ƕD=Iï��`��8�j�,+w��ϱ�ܽ�ѦP�*nrCY4�H#ʈ���`:n����S�˷=��jK�:1U
�6o��&	��9�
k^�����Yp�s�r�44Α+���������{��-;�B;���N^�ō DZC�$OL��)@�f�T�&�1�G3*����֬��#Q�3�N�����q$}��n|����`����+�U\�!ML2.ýƟ ��>��>>�dok�.ʲ�3�V-*Rд�&�pDr.(��fʢ`�fq󥶣�~8��/�ʛ{.��_�=�:��u�TB���G'��<{ic�:]�:�j;��^������?R���`J+��Kÿh���;=t���&prjLKʝ�nISi�/�=l�tH*�7�y�R�Ѥ�tP��o���ؐ	x@�E�9!L���3K�z�qz��X���b�+��Ɓ�)fK��B�gR����;_��0@�j�R�9q&	��zWO��jE���;Ja)�}�b:	��!=��9V;X��nG�ZdS3N�;�㰂"�cq�������r���@���X���۩�<=n�9T���9�[l�VC\��5�����~��h�ף�����Ǭ��ҢD�T�.;�A����=`_��w��:vyF�J���`TD�x�{� �LE���ƪ���	������j�E[�����d���8�g ��s�9^��u��5Z��N0p�6�4ƶ�𐜛�*M'=/��h1�}@�/��)�G�,�7I���dA=�) T%�gdRHk*b_�����h��U��P��8p���/��Q����׸�<�E�ɿ`+��<��[���N��*g��/=0~
?<�5P��c<ycI�����d4{�� ��/��BD݊J@G)�j_�̆��c�A�@�&6���`�h=q��G8X9:J��
C��J�'�6���٧S��5K���-<��$�ʙ	��-ZT�V��9��h5���o��!S�$�Aa�Y�L #���i�\<fzf�L�kV�ߩ��=�&>oc7��������M�g0d��OCe�L{��.Ϝ�}�+̅��f(�<UX� v��r�PC��x���,���S�.o������=<��40Ű:��[�fmv��nf��"���bI��LW�K���De�ߵ'5whf]�����K�b�/����q�}A쫂`dI!���r7 C�G�+[A�Vjz��U�]7S%�BJ�營��"SFZeTu���ECo�*ݼ�n�