��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��VB�#q�@�;<t��:�[-���&��5/(���{���i�9�о=�%}�~BW.p~+`�l�`��c�����eB0���iأ��䧽�|��b��`V�C���<9Bʥ�_,̣�5\܈\�#��W�2\ ��S�`g$�1�بN�=�W�y���_?�(4�R���Uܾ"P|��S��v��^!]*m^�"��@"�K��&�>2�n�h��kAŬ?=�1��X&m��R�Ȼ@�b
�S�J��߮{6V�U�5��SD�D���mc�$������)��ÙAD�����z �����W����ĸ�)���~!�^BJ�\VsQ�G귂�	�8��a�X����}������ ����y�a�j�M��5N�ym�t�g=�k�ի� �¶\;���|Aj��+�!�6��3uf��sV(�>I*��q�����E�7�A��ż��٬�'ƔM��΅;�HU��!=��T���@�ZRs�Ȫ	4�Y�
9ۡWlX�C�2N!-u�H-NY%�GË����<�;�J�Z���ϑ���'S����b����h@��n��B�;~2�C�n������~V���Z�_�ݜG�޺���� �&�<b��Fi-�?s��p'ʼx�
EߐS � �ai���iՏ�Ug�@�f��G��J�c���?���A��E�󌅟$s�KF�}]�������6�C�F^��cQ)�o�k|4xT�@k��!�|�M���~FNV�UoY��P�/MsQ$i�6�	_�:p�^���$�@u�K�y�/X�h���tَ9�
O�L���sn�_x�!������r TN��㗭'�H���v�qs�_�X�J��s�uV���=ڈ0�9��8$��לeL�+�'�����M��S��%'���}CP|:��>�#��g��3� �h���o%�G�A��=*<.������?�-�#s
�𣰷&��w��c����y���y@��
R��]\�����	m@t�b�:����L�C���h��������o��}���o��'����a�p5�G�i���"�hww[f�}�����ȴ��t�`:�E�1:[�
*-�w��f�E�(� �?k���A��\� o�'*LX��DH=�.�ejбߴU}����VdR��s�����vx���/F�]Z�'������ |��[�ɻ9��;�rGҮl���P=��[�'3���!�faδPe�;<Ix��� �gYs*�Xa�x��.V�Q|H�?u�Cc\�TC#��l�g
�Βʣ��!la9e%��(�q��N�]$+�L{�OԆ�����z��4��ʗh�aq�̯�C��|y7����oxD�}�7y�c/O���z����_c����ץ�,����:i(|9 |[�TW'j��ɝ�l9Z�����B�k����3	��)���@
���Q&��ߊ��z�t��o�5ŗ��'��1}m�~�]��|��tL�Pn��G�.N�3�(�����؉B����A��S*�yk6I�iz��v�\䀮`z|�ϳg�LO*�]�ρ�o�z��H)�}OU�e�Hʣ���|Y�&ኄ�^J�ƏI(�y�c@8�.�'�¸���h��Y�|��?�]i�xSS`y? [�G��\���N���6�>6×Y�2}2��?�獜�G�b�	��(g�6�����#3��y�ɩH�4���?c0�`u�������f\�y�[׸I�H\٬
�!�y~�������@`��Ϣ���;,|��d"��T��|������6�Qp�Pz��/���d�jOr���[فKHD�*�{b���\�[�mCfrg��pвb6�_9,ZO��4�Ƴ�1���۔jw�rE����saW�w<�O�4;�EO��I�G8�T����:����FG�-��F�խSG
�A�Џ�wb�6,�$�����(���%g�+:��O��ѹ�9>��ϥ���/e�v��ʈT�j��j��q�IL����L��l���F�n�	߆kA�=��~Zp5'��Ql�Uɭ���'~��lA�� T��V�-0` ܀���յ�NA�I��1�0N�+�N�< Ih�����v�hZ
����'��}��J�Cɱ��1>?�QB2VQ�$��<�h�6�J����v1��/�W���$ᙕ���@Яv�M��T H�<�s� $��Z�g\ruw��g<_��J�:�R7�^Z����{�,!j�o0�s��[v]u[1��'](�i2�r�]_���rnֆ�~��п?>$sU�J	�i����\$�hWP\���ns0@���Q�H�%p�+�&T\'����y��ykHwݾD
M����֝4�v2�P��YQ�2�N��i� ��F��4is�QHڼ|�������:��Z{x2��$8����x��B��ғ�n�K�^�AZ�ƌ�̽M��v�&�(.c��S5@.t�|�9g�i��*�!��,��L��r�9L�&t,%e�1P�^D	m4%\l������@��$��'�ȅ�͔���LIcijis��9��C��I�*Y�<b:)E]��K��Z�S��ё�}n�U��M�{-0f�sm�##�WQ�	�I�ol������xEv�1�k��d(,�$kG��"�K���%f5�z��_�� �xK���o���6c���iH+��H󞝤p	�����q=(�M$�p��'s�;qMY�F�s1�V�ұ���i�E~m�&^�-`
�t�fs�ܜXDb����%e}F>&�ڳg�����
�=�P�gF}�H���f����mŧ����5�f�s��R�"����c�B 9�ߠ�Kp���ꇰŕI�r�p� *��to'i �۷�M��P�E�hF��G�B�*���/�����F���l�8����OY�ѕF��)���� 6��NuW`6��3>V2��c�f`�.��}W�9H��V����������A%��L�%�}���(���K̬I2f<}���OX������!z����d��	��JrW5