��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȌu�(:�b��%[��$~�c�;+��~�AB(�DΞkv.�_�O������&��x�w�����^܋��U�dUjȫ�j��q5�#~9�w	��2�qt)�'��svk�f�H�>^?�Ϡ�S�����'#v������O���l��G�0?���.�t���z��NP�jTH�� íǘ�n�[W�LEi�(���o�G��)�\q6�<p%f��+7���M�G�c�ƀ����]�~�J���M�����9�`�<dM�\�r�~Z_p,�����
?�~izP�_���'#�x���H���鱠��6��#�%QX-��?�u_��|�pa7����yX��q��ަP	L��o��r�����Bp0��$���z�Gɿ���q����/��i�Kd��]ڿ���*aw>Rԁ���C{[�hm�_F<w��r'�R�&|q$���^��{��W*	��e�sjS%Wt	����Oc�@4�D�1�::AR��P[:CIG�h�{\��K ���͆Y-ӧ>x���MB��N�"��5�ؿ��H����I�}�7�����U#���X��=���ߏ���_�<n
�o�t;8z��^�gw\318L�2%��9?+
Òd�
�t7n�sب�}�+�]��OZ�m7ө[�,�^�~L0��@_,����dQq�U�<!�m�Z�:�G�� ��v��i-�p����c�տ�#�b�N	ơj����P}#� ���ύ�BD�D&�/�4Ͻ�M�݇����H��4�3�}��.�������<a�QH�x b��@�%dWS�4�7�ye?bfl�`���!e�� ��/�c���~��'W���,]�^o�_���C��j6gEV뇢j��cD�f�
��Py�vE�c�g��� ;�f<��-��Qm	ڌ��i��~��ay�o�t0�l�|�f8h5Y��m��U�_�^d[�H��g����a[��6�B�����"��j)o9]_��GrU� ��/>�c^�y.�Fg���Q�0��N�-�.�����O��v�b'%�>-z��Y�+�{�(�����0�DC�� J>�%����,���]ܳ��(�&�{�sl��-G��p����<���N��2QF�H�,�;2S��J����۸������Dbh�P�X1�c��C��N�<bp�ࣄ+$�0���Q��t;+%)���C���'ο8�C��������b*�D ��t���e��Q�Lu�%V_ȿ؍�c�Wt!��ӭ�=�j]�˹���������r��܁Ifv
iUCU��/�z��^�U�rMgN9�(�J�y0���fy�K�\9��{�ʼۘ�cC=�U�;hn���Q@�\DX�����I�x$><��xz�u�Ǵ3�q��j�&z��2h��D��D\�p�8Ԭ���䭧���	E}OK,2���1�(�R�X2�/�DR�
lv�z�n#�:%g�2����:����2��E����k�c�S��`W2SL�VrQ'�p��pWy�j2'�}�!H��x�Fn-h���%	Hd3!�W�dj�zFs3��>�"�؝��:U)g6�g<�d�7h7��L�tJ����oH�]Pxӆ/�"�	`7�������r��3�D��Ėm����n�	M���ƈ�\	�9�	4��r�+��'�w5�`˹^��5��e"
Tb�	��];�߯0�7k>���Q�!���~M�a~O�����)c�0�0#��\��5l�0ԯ�r���i�4�K�g]6��U �?p���TT�s�b�u���L��2�F���uW�d��b7݊7��2ț���c9^�\�T�\B(
�ivU˵9vpƲNlO�]�y�����k�aS���]^ rtv���� �t�o���J� �U�^����m�_p���ټ��H��&���{���U�2���sW&W���BF�{�W~`��l۞�!�ˍ%�k�.��q�UӻZ��y�����a�3��}'1�h��ttl��QDnrl�&��@�9\#�=��Ǌ�I�n�",� ���b<(49�u��L�Ó�J��@�P��2D�0i�:��Y��^Υ/����k����9��׆�SB���Ӭ_1Eoz6��v�3�阹�o�jf�;��I,���L����Fh�kq���C�#o��� �6�œ��^��%	$޼b���";X�듕�|���wx<P�iv�ͬ`�$j����e�T��R@�� W�_����;0I:�^�;��H��߸�5T�T$����|l.��*����q��g�$`�7G�5zssN�B�8�,�C�K�*���C��R"N��]�R�v�/;6��.��F��0�U��޳oS��XP5���E��mQ?�~�]�� m�� ��#�9���S��������h��<�|�I)=�d9����pP`�4���".���0�|��O9��Vkvc-�����iz������f$��$95�����PC侬>�����u�d�A4aɀ{XESi��A������X�z��ґ��t��1�b,�|�g{��6��H���\S�e����{�������pg
`�H�UX������*�c+��BŸQG)��m�]�&|Q�\��8X��_c�Vu~\�\9h��R��olϑ.�=I���8c�n�l���?�^W$�@��O��nO؉'��`�o�TţX��������4�tυ�2f�	*�����e�>=w��/v��6������P&n���!b6�#������Q�"FJ��s�l(�M�-饱xG��L�oxZ�t����jap!5N��_;�Y-�"�����H�/���D��#������!'�m�W�kZƕ�7O�p�jŸ"Q�m�nԠ�H�1�#�"��d���G��v���\���0<<qX��.E�ߦ��v!;5h���d@�A���r-�og���q*���_��	��@���n�!�+�)���,���<�
��Ls����I���|��k�W�C%3�|4_]�<�hfA����6�eL,�LIŖ��@�^���N��kl%�y��:�Un��ߤ�v��UME�
h�)���y����,{S�z6�2��G��Ǔ������ݡ���hW�ҷݧ�H�ȉVԴBA�oq
6������v5����RzC:�ύu��k�d�3��a�?	�1���o ��`�|�[:[ˏv=y��k�s�bagy��ܴ�-�����?e��6�fJƪ�q��:dd�DX�� ���N$;��������?�0���\�^��ط�\��u�9a��*��j=d	O�p�F)�=�`OfMۀ�3<��X�K��6���m����T��qܻe���sB��U)�v�F��́���	��{�d� ��lu9���6i��b���<�+}ߗ)]��-cr˿@�ӥ�X���<�k6ej�����2W�i�-�5�g'S����_&�Q_q�#%�r�N� q~�v����e����@g��f'��4_�q�������ͯ�����	PӲ�ۘ ��l���cʣ=�(F�wv��ó�y��!�VH�����j @�(�uC�'�"L	 �D�vMm�Y�/0󿬰����.��?�"�Z�D7m%����Q�XZV׶�^	ޑ�y!P�3�~���N��,�z��[��Ήl���,�=|��������\bM���GkL��"�u�wSe��G��o��2?�Hw��������2�VNj!����~���B��a��e��+�h�f{��HC̱;�����6��|���>#Z��8�[E��h�vک3;@������jyw�⛵�1��ȻJR#U����o]��\"֏1=�c$E3쑛�{ҡ(mG��*��D��~�k�r@4�'d�y������8X�XRgsq1����*�XBAL=�`�IKG,ۣ�|�r���!5݄��X� B�P>l� DOO�ڇ�٠��7B�F������Wb�����c'�P��`;3�E8h�y�K�M��L��˴ �T��=�F�,+Q���^Eʝ��_4n
�`Cgl�vCԠ`�ǭ��{�38��d��GM,��[c0ᄕM}
w���2y���7�1���iL�ϥD���u^�} /ysW�{��{�l����k�Ǣ��(���[W$My"r/�x�3�3hD�[]K>%�)5�����m��Z�T��5#����;�a*���U*ߓ>6M��'r�3>�����1-N�dnc�%�Ms���8�˸6w���C3�d�~JO��I�~��Y�Υ4u��T�s"�CC�q#Y*93s� @��������� '1p S���A4b!o��Dŕ h��@+\���e��\��_ ���/U���P��\� p�\��rV`!O�����5��#5�C"�<��rbpU61�o��८)�3�7>��'�K�_���S��v��
t��C۠�g�{��f�7P]���o�m`��oƷ�"z˻��Y����,W�nD�=�"�7͟�c+CP�p������Ga//S`���s+lA��6��]	M��7�h�.g;-�_��`�`K�B3�.�$]��.��� D��]k��O��Ќ9V��ޱ���AĚ�p�Sӣ��*'�$�i�;�Xڹ����$�r�i�m�88�����.�!���>B5����?6Hpbd��*8��d��(��"B���m��<��2�m��4��y�G�NK@m��鉦������:�X�F���x���	.KB�-1��K�M�x�(V��/ tޡ��Ȇ�u�8��A̼��!��-�2�z�Άh���a��ڭG�M�b���E�L�(���q ?�23��XݖiX0mrʈ'�i�(Mp(��ډ��U��N��P�$�A`��h��|=s�B�2���N�#]4�>�W6)i�������0@��ϕE輧��?�Q��V�������?�ɂ��@сA��UA9��܀����dJd;��B<iI,��7�ǀ�?�>���Z��\�
h���P�0B	��#���=pV<��7�ѠWp�L$"3�)�b���+-+�Y�:��èY'�������W��t0�gǽS�+�B�JK��徿{-h�w���h1 P^`i��m���e�?R	S#���G/Y0����x�1�q��X�8c��e������[}�g�<���!����C?:��z8�=���Q�#���*�͘5
x1$���֣{�?�5C�U	�kd�����}�U_=M�O��[ȅ>8�6�PzW�Rچ'Dx�k�2Ԑ�|�����x��c�r.@�'(��Gh��G���{�o���\�����o��!��ǁ��$5O���ͧx��pO[�\�2y)i��X�4�#�qnbFA�v��\�N�h���L]�g`��.'s�Ch���	�.Pl.C��֤�2�� �68��"�vQ�\bsE%�bH�?�&�6�qE�G&%w������n92�QsM	捧 F��z��`|~�ISKM���)�-���^>D�����o���%�Q��l&�0c���A0�@M%MĬ���+L�}Tè����x�U����T��;z�u�[\	�}ys��73�y���<n�<���@��@�q�#/
�2F#i$����J]�j�Z�$���]�m��2��s֛;$�n��g�
SI�E|���j��p]�վxz��8�4]�T�j$�4��i����������TfeB�;X��H���ŵ�,�[�*��~3Y��@C�?v�iEWk�f���{��p;���
�.F�[�@��9����r�Ò�zԼdD3L��p}PV��<�5�vC4�?�iB)�W�S�΅R~m1(�;g�Dr�ϱv���[ב���E1���am�ꏿZ��h���>���C�R�=���鈭ʹ���������[���[�\������u������"���:��u �ׂ�����bi0?AM���Z¯�`�����O5,m�3D�'3y�K)7�?���`���� �,+x~��<"Ł�\�a��1����֍J(m�^������LK�t��V��r����}� �Ӳ#��Q��&��̜&��AX߮Y^���r�x3)�n�-�O�4��=ޯV�Z��*�Z3'
"8�Lx�S����i a��𚿚`)�@H����#{�qw+��O�w�s��*-�����TAN���h�,�>*>ف����bƨzq�!��)Ȋ�Pג廵-���j�����>���A��ǽ�b^��J0#Ց:����?� D>����D���ش��s�ɷ���|Z��;�<����r]��(��+^&mW�9b'ǚ����ϩ��y	���������vĊ�qP�9W7��e����DZZ���{<���C2](w*���O��ׄ�a��b�&:���n.�V�[ZWY�iI�i�N�gl�,�`h����^!6p���K�(�/<�����jH��ƼD>0���m
0�Q�yE4Zn�PGa/�ݍk�I(�� �V���o��>��^O��8�4]�B�Z\���K겣ki�>{ѯK��ntW�mw㩾	1`E��4Z�Ǭ���LW�"�8mP���Nt*o:��:[�+Ѭ�*��Y��ǫخ��䳀���N[�{*���O�:��p�.��w�[�܅׬�
�qI�Hi��r��|����DcI�~p�\�|��P��u�mv�n�o�����
��������X��F�|O����g7��?OO�߂���t
4�xA�i��y9��(*iX��B�N��ITD�=��T��H,��sm�ė巏`V��Ȩ���բg�MEC�&�k�4� "�ޗ0��¯�A��	��nF2�_3���'��pnD�g�����؟��7b�BBʨ�+I������������m9m�%���'��m�TC8�m�b�N�8G�ٽ8��b*-C�.��6��UTr��c`��y��n�Ub,X�#�Վ�Ċ��H�����`':)���OL�a�5�5:�������
�����.O��l`�kF�/�����0{	�^jRk=)iE��g������$�r���T��.«��n,2��y� y
�9��(c���g&XJ�!ڡ��f�̎�V����dmG���B���whs@�cH|e'���;2�_:���KPXF�23_��7���6�4GM&;�l�*����j9�I�,0l���x�Q��C$XHC�0�M~�w��%!2K޿�vڏ</��eh���X�j�c���������v�0��$|���GB��o�&}_�.��w ��l�|�5ȷ_T�w��I6��3ݬ��<0�3�`���Af/�u��J-�}�W���Ks8����j��W�Sw"jO�C��j�L�w@�ɘ���`w��`�O�������q��v�N�J��B�F���E�E��+p�H7��j�˹~-�$b����,mVF�+*�p��z!-Nh��*�"Gd�ф50�����H�j���+*��`m���A�:�r�*���z�S��12C�=�aX���uT�9��绂��xvqծ �S n� �� �Z��'�;�Hx��>��j0�ƻ>��)|H��yY����`��0V�9����҃��^?)#���`0�(f�O�m�`B�l�|B��M/���
�L�,/����="�Q�(P�u;�z��q�⯽9�x�V%O�k&ĂGM�cC�FSd��>k��[	(Y����y����Z�d~��&׶��V1\��n�ҭ��P��Vu3h�C�����a6^�1�ʓ�}1�B���t/��~o	����<E� ����Z&���8��	lGY_��gά����r<�<�e�O�ծ4���gD�+��6�~�¼��NWX���Pe(E�["��	^F���֠lpM�c+U(���
2�M�H��-�NZU��B{�<̡����'�,?i�TS�c��`���i�K�J��s��cI�H�Z�1Ɔ�S�S���5��m8A��V���=^6p��/���?	�T���a���9j�Tټ�;"5O�>
����_���X�����[@��&v(����lQ�O��t�����r�!?���Хjg���Ƿ�.�]�nnO�$���!t�@߹��b=��s^z^����:���2����gkKx���Ȉ��� scb	|�tm�v�H��`[ѹ�>&�(������%��XM��#ϸ��VI�u~o� @,Wǻ�aU����(:�w[`����g��B�w�{�����jS��.f9qP�b��0��?C�_E3o�5�q �e���Ö�RG#Q��� ��Srx���\f[����5H��ľ��y�!ނ����/j�>v�V:R+�u�_Xܿw�$Uo'��aډ��������3I�I�)���F"����8��̾�i�e�<O'��rv$��;��`�"�S,FcϮ���}���!�⏪Y��/���g��IAJUG���!}+��Y��n�՗z=)�ÝxVI.M^�ۈ�R�Q%Q�F2�'�$���'+�b9���Fk�9ad>ۿ
F]BXGH��8X�PC��0��Ίl��ۡ�k��f[���f:(����1"n?���H����i/;�5�Q���f��v(S����w��2_��W�#��y!Թ�/�������L������3�aV�{��z>�����ql�F8E��%���@� ��y�-�LڞC;dz��q�C!#�SǤ��r%�+z��XN��CК��"4�]�l�&���FT��MH���JMs"�8�3&8m}ֿ髅Pn��Z���*i�� �xUm���U9"wʶt[�� �՛V�>s��,jʬr��P�KQ��V��:� :��(\�/�(b|�}k����[�n;��qƍ����'H{�H&R�e�.sN��b�X�V�'w$���4��W��s�QX���W5C��ΣT&�~
�G�왵���b[]�a4m�6����8fj�ͩθ6��3����:t�n�/KzT�":�]T��čE% ����U��	�|><0��6S�"�2H�^�����#�b��]���a���`8|����$�����-Y=��DD�ޱ�����|6S\aZ�4�γ�J��I���֋�κ���`r�&�U`2���u�V�;&�#�A&�r�@�w����Q��'c{����j�f� d�P+6��ѧNL���-1����Q��M�Q297�l�Fs��T@	TbF	��Y�G�~�rB���m�J	�rC�j\��ռ.�����Y�����%G@O�x�Xxr!{^O󥫽��<�]p'�QBt��3v��ί����\0���3���ݞc#��ᅦ`K&U	#l(� ,������%e��d?� �R��c��p8��y[q_��M���O*ڹPN~a`}�i�+��w���Ta8U�9퓐*�lC�E7h�o�{�$��]�aȶ��������s�t`p�|v�=+�9��qP��$T|ޚR�"�y�R�O��/��7�r���t�.�sы���A�u��v؋!a�{��Yy�K�}#���O� �p��ql��G"�˼��@	����MG���>��y�*P�fc�U���Wչ���W�Q�;g��]�	+��&p�n�9��Wj	���P���+�9����Қ�;�x��K
����4<^�~��w�A��y���C�$$�&T��L�c���u��P�Qtm	ب��� @����uK�7�'��GZ��i��7 b���%�z�������5p�D����!,�� 5���:g��ǵ׋�Y`��4������-Y�A2w�Tz��hzs6u�F�'�Z�5Bپ�i��?v-���Y�W$M4f2/-�y˗�V�X���a��0����m|�<���s�jE�8g�J�I�#6�{0�p�!�ߣ�M�-Jه�#�͹����������C���)6i��v�aࣞX�aW�M���yq���٨C�6�̻�r��o0���k�о�����м���4��r�{'խ��!�	-����=.�~=�H����}���x-a�_���H�|4�d���#Y�K�;?��
��h���s.S�[���l��I��h�3"��( �Fe��F+�5��x��pO%�-ir`N��q������m�v��.�G�W��Q?I��_��i��X�V����lTP���pJSf���^�R+��|W�*���o7FAq�E�O����+�g6�-~�	����T�,�:��B�c�[����,;�zܡ��AA���C��y#�#�ʾ\K�g����m�^�����vF�hR�S�����ii|:���S3�&���I���Ey; ���s�R�g�H큉d2�[	���d2al4���x*�i�p�~�8o�~\��WBF)b-��K
�a��+��8�J�ZMg�^8P� )&�mr��G9vC��%�a�
��׷zw�S��J�E���Ks���<�=��S�;Qӕ����xK��T��>0�}��R���R`o)V��"�s�p֝9CF�&:���$��=$�b��!��a�XA���y_�nͨ�������;:k�7�9��.,�d�����1C.�.���.B.�p�26�:�����!ί�fn�X�����@(W������@NwhQ�3�{x,*$Ք��|O^��`B�G ��'[иE�~���pO I�SPr��}g�i
d|*��0o�r5|=[���.��}]�x��҉��0�K�n���%�(��r."��ݯv<erW�,P��~���n���1���U�IF�>��WAT��p�U��{�zK<f���Iƿ�$���1�����(n�i=�k�K�xv�M%y{2���9�u@��)�T��y��Nޝ�:�_�Ӟ"�>��x�w�|��jf��,�]Q��d�ER����Lj>��S�?��ǩ��4��4�,2_�@��ؓ�{M��7���������wWnќ�=U+٢��W+�����L��7����K0b���&اY�Í�Ȇ�\�Ȧ�mPS�Ƹo PӖ����BUVF��S�i!�)�j�7���4�Dֻ�<��B���j�_h�ɐ�}Dç�0�L�!$;X�7=
�����I��T�m�S��U �Mą�9@a�(���K)�r��_W�(��.o��JDl�!��}�&ȐZ�0��0ǉ��ʑE�P�0f,�f�G��i	�k\n|�R�<�4����G3����`�*�ՎX[K�mQ�f�7�I	�m�EP/�`>N�p�4T�)F0u�������L������>3�~
V���K��y[�/a'6=]3Eq�;V�e`���PJ,ͪ�|�?dgz�]2<�����Lq���������{�zB�U����c
�抨������'�:(9�P��@o�ϩ��W���$ С��� ���h%ީ4vJ��,�T�]�P))/օ�����!MD��'���49@A����F8��z7'�A�窅��q�˒LI��sMߨ� "���Y���v����mC�\�Rj��0pY᏶6(����eJW�=��1�����fɋ�ǅp2�?Zg�b@��� ��5	�,��ZZ{�r[n�rv�"Q���ᘲUeA��)� 񁆟��/ǆmR�B�>��5]�B(Tf~$��hC�!��Ѹ���A|-��
�\[�0T;�J�� 1�el�1i7�y�k�yi���!���*�l��w6�$rV�q��7Z�>�j�/�w�������ŏ�|��`�j��n�i������<��G��z�-�c<���t��M�~(�z+�Q�۰-�c�
�Tև�|��Yн	��+$��� ~�J�����B��|�RZ,�����t��Cv��ۜ�tw�����	x	�Q�9�=v|����~�N�1|��)9��mTB��������׭�0�V��_��LA��o�*6h"��=�&u���b���"g+�e'~�C��L�9"��g���:�$���;��m���;F��Th���]�G�S�AG(h��8I��O��`� ˔*����W��={�W����?唗�3�P��� ��8Q��d���};KK��\�I�p���W}DZ`!�a�گY�VɣV�HN���֞�E���g�L�;��J������ͼ���7Ysl?�����ͭ�����ϷL����	E��f\����Wa&B���n�����~W[H��$�e�V317 *W�[p�����C�*��_�.��/)w�Q?�$o�M�H=�J�b8��v�V�
����H�)��y%N~��������W�wI��&���}�9�,�	f]n���q?04�
��H�����Mm�=��]��-������X���glNM�@r��3t�$2g,�0'�L���R
��J_Q��#l���Љ���Э�m3G7`�U)>����3��_�����7�L2m�K�J�jh�>1���(�S���#�����Z�^�f�''��P+��,:ұ�D7������f��_�TZ�2��~��د�o�޷+��Oۻ���C��k���>��(�bR�T4sI��=&!+��O�@�y<�[�J}8*���W�B'0!����S�t��MM�'�� �G��R�t{��TJ'n�CM�-T���R�&=.{����H���W�u��6��͢'�+V�~�K�H
oi�sܑe��bz�����֡�A�p�p�*��P?�,$go�����3du	F�X �I<�]��HP�u��O�b��ّ��%���u����y�f�}z	{J�u<�|̵G& ���
���� <��/��X��Pع�����P_��q�(���/@7ѣ�Z�ݚn_Z�(�G9+(ҿN�AԳsP��Ms]q	bf���۠�QK����^Kq0��+[�H;�=�[�j����Z��s̲K'�����4'ϟgC>>zW��T��I9�Ou���u]k��a﬿�A�c�q��J֝�c� �PU�]W��C V:#^T��;����"��\����p�{��A�� dd˄?�g1Vƛ�y��}lJ;M�V��;N��Ơ��ŷdL����I�,�Qo���"��u��9Wy�	L�!��9at�Co���d�Z~�aM�j�z�� &����t�iL��)ZCg��zvA�9��2��|��ߓ�&���$\k4
��]������C�6��}d ^(�;*�^���yR�*%D�j�r�۞$؞��R���ن�|��fK J�/ۭ��ǆ��[zx�8:�x�t�R��w��g�
�E��ʼ��rD��F�VcJ>�A;��z���H8�ܐgF͈!�����3�P"�^~-���`�������B�Dz��;��,��E]��n�-	�?��Z���U\����E���Q��ⰤRpRQ�ƤLcTo��/�{1�6��a8y�>���؝1#O���Q5𷵡C�/n&��B#�[����Ŵ��0�ʱ��pj�`�K�(�%%(��Hx�T+����0W�֟Vs�@gEp`��=)�y���
������fR�-H��C���w-��oh��ٸ�8�ɂ뤘��Dt�z��G5;�s�Z�hX���vyc�W���s�����Q�4�҇7��(^���ή.տ�q��p�����4j�Z����f�f^3Nm�|�ކ�=��4��-�i-�­��]t�ڸG�W�������V�]��
1���p���9���U�}��3�Ɩ�"���$h� 9_&cO���:#��Y O�����"'N�磫.�e��aL�`�@G�5WB1����b]��T{Ju�[q�I�:�N?[���e3���~Q��r >�0�M����iܴîAo3�&l�g��K�0��t'%�C�i̳��ԮtB�(��@�*a����Q^��x�*LR{��`��5!8?g����~�@���}h *��ڙ �x�!�5�B�?c0��:>���떯���sѝ0��s�k��"қ5�	\�/�����J&�Q{�U������<!�M�H.8�b9�y�rGާ�x����u\�b6�̕�@Ɵ��'$�I�_�@L.�����%R�Y`�hZr���R�vn��=[�	�*T���A��xn9�;X�r6�Ewv�3t�춏�1��?]�9�xl뼜;o��;Qz¯8�s��¹oO��(S��(92�J�.��� �i(֠�\ҿJx����ޫa��J7ŵ�h�?��h�Xr	�m*�����m?�k�,���8�j�.���5����Q�3�6�,������x�������4t0tE��NB'<����mg��b�]��W[���g~e�Or��As����_�L����
�
^X�<�<xX����[H��D��QT*WE����7դ�*���$�Ц�n;n��J���:�Q���)dm'c�g�א
��y)��f	���_��k���,���O�ô|��}P L��*,��yo�E����#����0��OX�M�y;긶�E0,��#�_`J�XY�K���U����Z�
0O ܓ�|`u�-�+Y���%��g��5�����;"m�m �����B�g$5J����<䄔���|�	��!Lb�\�+�?#E����R��2Q��\��E�\��D�S��Zj��ƎޘK��sɉ]{]��'F�S�7vSmD2�We�*e�²�9�A x��ߖM)Sq/�B�<��8�3o
}��fd�2�-�:d@��J$�ڊ���
�s2-���1�k�"h�op�l�z6ﵞ�Ѳ@H'���/�u[C+g��/+�7�f���@�8�Yص/���eѴt��-��0 E.$E� �RF�㴴�D'>9��e��v�����{@��`�q�X�M<U�e.|��9��Ӥ�Wi�s�H�밣��%��4!:��4A�y�}����	^�-��m���+��M��H���&d��`�Q�SU�6��{��#��oќ��.f�/�w�V�Co-��^��R0 ǒ�5�a��p+{�,��z٧��C�5�����5�o����u�V�1��w�Us,}$�.ت[���	�o�1!��b��w�'���Z/��G��1~Ո������'�$����������gr�� �nf�����#�6uءn�~��$���jC��ɋ�=_��G�:�.�ߏ����`9{�����MJ���m�`|�E�uO��`�}�H7V%��<�Fɸ�.B�4O9�����y��_8��}�ed��,���-�&7���>E�K����A�r�Y�.>�̓n�����y~���KT֋��CZ�w���\�KO�Ѝ�v;V陫�}��Q$j�À]X��oi��!1iz2��sPv�9�=��Q��!0��lv�ϟOP�m��6��|���^{s�XG/ؑ_���f�|q���T�A��w�/,u���x��Cl��P&��{	�c�{��0�w��'ܙw�H�EĚ��r�5��5y��/d=!�
��{:��I��CBK���?�ޝz4T1�^�:8�%~�oKk�+)}� ��2��?����1M�x�7[�䇉��N���a7�Ђ�E^��pVT:��W�d�:��󔌬u��.Hn>��պ���v4�n��.0uh�0�VS������9U��"�d�Y��K��aW4>|���طj �	Uǐ׉�%Xr
�F�TEs�EW)	�xM���0�_3��؜���u���h�X�����O*c	��U��$<>��4%I,�LH��dgc,�>��X��m
":��&Vl����_`�Zh�A���Z������/L9~�	@}bY��d�D������6��'��5�L2�`���3���G���h �ث�Vmd���!�M��dTQq�U%������C����*'��<� ���j�!�� aN�:�k�Tpҭ����>f��+&egbXq����`ʘ^Mj�{��B�������@D�گf!0!����Cz��|-�m�]�b}����-�BL�V"�c�����a�V�H�QE/1\|��H��}S��,j<9NR��?t������/C�\��:�	��U�GIM���BNb�g8�5)h�mڪzh�4��V�yY@�A�[_�[cO�a/�=��ϋ�$֙Z�Ć��
�N��x�=B�X��.���)�eT/n���/wG`r���+nS�Ȁ�8�2�*ټ%9��ܪaP"�KQ�� ��2��׈T� �[�{�. �	Ba���X���9+��X8����p�o*yAU}*��<����>e��?��S�46杜{X2�`�&�3�7X��gD�?i8r<e���;����X����S���@`{�i2]M�)��{j,R��;���_|E7 ~�!����-���E�a��l/QV�����SN^��A�|�&%L�.?` �U%7�����C�Y/��	+a|4��|mp���&φX�r�9���N���!Z��_"��ȉ~�[\i$�:�q�N���a[g��_7�~n�\�̿h>N�eǸ�q[Q��B��o�``s�`��w�әH�z�*�ֳ�C�,=��Y���X�ٷG1�)�?2�kd?�^��Ġ��̅HO8�~V�GX>h�;+����g�n3jI�h�9Q����6�'�j���^���{s����N�Wsv�U�8
��:�΢d�(��@"�mX��|��?�Z1�|���tDb����x���T>�b�ζ�L�8�Y�/0Hfo����@�㧱����hv�U�{I�7B�Vf^El���rnS�2,,�*懠��w�b0U�aq'(��5k���$������M�}+�@K8���NR��� ���9�d��uհv�lu�Շi��cB�<�ȹ�z�!�_.�g����ي1p0�[�4�Ei#s�`�CA�l��Mm+*��$V
 ��|�^�+8G�.�{��D�Qj�&r+$�vj��T<�g��I�w��ǹ�ل����]��U*l}�������Jc����J#��߽�!�8��M�R���/C��j��oW���A�{���KQ�0����q�6X���]�k|���5w�Ib{3+{(D�Or.��-��O�K�I��X�{��R<&�~ޫ��6/�ڇ
�NR?_h��~�DN�+1�`�`!�굈��[m�+$B<ފ�������,�'��F��&E�I�-���4}�F�<�`V ~��L�eF؜-%5�����ցUr_H�Ȕ�1e�;
v�5��i±�Ro�|pN�[�i�@��ӓ��ytҢ8�&,U,�9�_�s��}�o�%��B-�gc�E�����YCY�C���|�&	=�C@RM�A?O#����^�9��]��߲p��.��ǋ�h��2jyIc^o����^�y��'�n1U��^n�0}E��J@��eJհ搂ʘ��/�LC���B�ʸ��&{��2۝G���a.����X�"���u�2 ~Z �L���A�+F{@���$^[�j}k��Y&ʂ�'��}CA�8�����#o��1Z�㈫�4����ܞ��\0��ET/ݝ��+c��w�(?@8��`�#�!BU�?-���4�W��	�g���)�x�>ga)�n��� ȹ �d��f%t�m�����iDC/�Fx
�r5|cn��sW��DX�A�{����*+��62T9 ����\�����\��J��BQ>�3�� v��^ۤ�ؤ؂�C���C�<�L��tظ]���:��A�w=�:��s^<V��%��T�\�b؋$��i�+����ښ.f�^�̷�L��H���I}c���Nb[�n]wL��0���>!�V�C����}Ŀ��^�|��h���D&����)�D+n-D��t[��?�}�d�/�.�K��/t#]���	"�^��_����[x���Fi�ڷ��u��qp�V�{�"�7�vj3�&�(M�d%-�w9$�\}��_�96?]� �\
3����"w��( j�kU\�ov�YMl�{��07FJ���?��o�w�,��+��u�Q2���C���E1ѕ��[5_�C����m���<��Wpx;�:��t���9y��d��`�� �b�/0�+N��c�	��j��wRۥJ6�N|�f_'�����0P��S�Y�M1����)k����͍q���Cڗ��zQ5S������%��*��wNO���p�,�D�_Vz�<�H�4���f,�f���Q�WQW����ϰҖ�B%J(P4=Ae̊����ey���r�t�;E�J%��n=0;�`�q�=�.�������+^�������ЁZ]�����2���Op�F�@¢���8��YD����W-NXI�8����ei���7��w�����:���M��4����V��tz��D,SXX�(�G����J5U��{��eM����`,�y��� �r?��k�6]|r4��\b3��`��xBt�����W�%�q�{t���D�q	{(�4��J�ˌ�$�]�n�n��nud����5խt̕�ydZ9N��	��-GF
�f,�pC�'�p����ɬ��ߔ��^Ɲ��(����M������RC��Yk�loˡ��C�6�$��Y��c"[%�,�f�%vDy?{�xeL���O�P`�T�U�y�#��乎Q��Y8��Q82o�T��l*��M�w��g���hɆJj8�W8�Y��{����O|�����i��K"U��@���Ϥ�����U�`'�"��Ǔm��������{�#`;t���2��I�x����/%�Q#eb.�+8]T��g��we�P�A���j`�o����{�e�U ���|��ҋ&������/e�)�ۄ�V�����"�R�z�;��~V���2Fh�P�2w�Ώ�����P<�ާ��wl/���)}��$�����/� ˺x�i���Zj���GY٪o�\�Xe'��|EQ���Y#T|�uTs;H�3�y܊�V1�\|ic�2k1�-n�l���|�,�����Q*̮x$w�s�䚭FS!����ޢo�Q<Z���Ք[#6/�V����p%U���;��K]FtU��w~9/%2���ׂ��6��փZ��Ѳq��Q5�zZ�h�P��"�

l�����u$^�~��s��F\�fxk(;�(��J̐���_���[�V���䲎{ezdA�K�`顰��Kc��D����u��	��E-?�a���Hȅ��Ѧ�PqZ[b%l��@dh�I�X��O]Ol���a���d�7�'T���`��ց�L�3�p�k����* �G�U�CV���P��r�X}J�K}6O�١s�(W�tw$� n��������%'��J�q&ADx�/���ܒ���!,��*0Y��0�YI�ټ>'>�ްO��=��ß#6]7��}�h#f.a؜���Y0l���V��[��X���na��3z�E��_���:�;%#P҃�s��W`s�؆��ՠ4�["�!S@rH}&�o�O�s��J:[
�(�/0�X����4��7�͠kGpg��q�������2�u�ڡ�Y�$��n�I�zl�� x��"�.������;�q �i�57O�D3x�hK��H�q0�A��·�j��Ҍ����]�G�h��# l�Q�;q��|��_(��QĀg�l��1�z�]v��I��]�
]�n����]҂�1���rD���\�
d����f0��I�!���.ȟ^�ȠB	.��eu�0�Gܯ���(�þV3����i�2��?��������D��d�9F-�d��`r�*�Ձ��Jc7���b.m!�� �yF̷fM< �J&��V���u�%���}�H\���R�N��+���������$��� o��y������8ɶ`e������k]���͐�X�n@��t�;�v���Sg�{2�Y}�di�>�}�'i�c�U��>�t�m���9ښ6��!��xkޤ�O��#���>����XG���5�A2R,����=q�:�U�U�ժ�����%ω>e�XNE�^!O	��3X�켪,�D��K"��RC����z�Pz�X,�VޞW`BKzdG,�b�k�R`[Q���?�Y.��a�/<&HA�
����o��+DC��,Nrs|	eiA9[��%�_���s;�W=�d��2B����<Fۼ���`(~z@�h�C*�b�x���f��+�h��G7�@��Z�N�e;!Y�<����>��H��:&<��=�Om�ĩ���o�
�s��Qy����޲�`�z�ҏT9������򪗡�V߶G>l�4��o���[U]¨D��.�zx�cŇ��:���u���t�(Q:�,y:FD�g�D�(!\���<�k5����i�"N��r��0A�uqȨ��H���X=���Y*��h��4��ܟ�e||�0��������Re̖��o�����2��;o���\���g��bD�6�|�J���ytiי��IbʙBM(92���}�Ǻ�����eP@p2�	� �2��:KS���x�J��z��U�g���u1��T)��7��h�?+�;(�B���Y:�!�K��}�!S�L���4C�Vz�[ rHlDA%F�]���$>�I�ː;VIhT�v����Q� �[��.�ڶ�,�Ҫ1ʽ�>sw��@��J�A�����V��Au#�d�ە.KѾ�i�/k}��F_���1OQ�Nװ��w�U ]��O�5�|]�tgٷ��˯�μ*2�X��p�Ocz:���}L �n�g)/6Jkh8�_/05Ry�ā�v����R��0P/K��,���Q2��"��=�ҥ��F��(e R�ڛ��5?o����h��a��C�uĚX��D8�����qbkր�#�h�2���9M���(H^ra�࿍9jL	���-g���wBQ����M��)l��S�~�~p��im��_����3+;N��MT�=l�|vc���ә��`+�]𞙃1_�N��L�U���B��\�����S����\�(Yeu�@�����Z�����U��{�}!F�~w�9�`48[�������擃������e+�bΑ���-i���b 2w�K���kt� ����U�ޠR���8�{�=sK�v'���3�is������b�ՌH�UJ̀W̭?�#���<�U��3��$gD �)M�q}����I�e����È7��T�^BHR��`����!�]���m�hשd�����A�!*x�L�!)D�t�yb`���F{�]��޸��L:�I(�6ZK�X��u�ꭢ	?�:��]�@e��i������
�����~e^b�G��^�E��EQ#�����/`�+��4��O��d"^'Q�/0]18�5�,�=�z"?���C�9 T�4xD�=O�8
�1/=X�$il�M��8{ ����Nj���oE��%2�
�S�m�W�G�p�
��Z��5i}h���h��{��f�����:�� P�����c�F΢Rv�m{�À̓��ўf�����o��-9S��tJ�T�`�h)����8[���`���X!�:�$�5�3,Vt�?�D�(Ϩ(�F����=�%a��R�p`��T�|ܿ�yJ1�lT!7G�+�D�5�֞��6��3�
�$A/}y�n5�_V�
�0�D�Kn|�+}�^1����G�����z=ɔ�5ri�?����a���X��zAМ��ς� �V=��Y�.6(x�6&Ne�0����F���AC&�4G:�9h�ۤ�8Dw{��%�5�z�Ո�}�h��]l��#��D$yM��V�<��Δz��jt�{E���2)�H���@z�g7�9)<*�S��Ne�M����˟A9�O� �M���^�E�O �7�{v�tn'���p��/�b_C#�n�9�c>�np d�ɠ����LB�7�s^�p~Q�j��m��_(1(���J|�^�32�+���Q���^-��؝���l��������d����+_���]^��F5'�s��XS`�;�'�<��P��V���y^=h��K���#��e��z	�h�T�I���6��l�h�_0͝;�P�ky��~�.U���q������'f����Ns�g?���Xg�7����j�Q]�߳��Pf�!�S_)�gx���읽a�v���z�#z�>��?�x����(n�X7V���E�%,�B��]tA��P���onw�8O�E���),B+ٕTC��+]�ղ' �̌"o�姏��F��jT��M��� �m\�MP''�e�d���R;�l��Ze��������w<�amǫ�� �c�3v��,,�Z���Ӝ�j�j�Ն��ko��1ה��tW�Z[�.Qڈۄ�0�p���� ~9Uc��<���oȥ�u� �Zơʛ�թH�%��kSG�{��GeL�r?��M��'����I��B��o=��V�2D��.��?�c�����?�uGʝaÍ���CH�O+LS��;s{����ؗWkF�����C�0��f_cz����y�<.{��._���/��zei��MPk�s���q�я�
�H��D���x�k�Xi��~d*9ʮ�~G��{�;%�^ۖ���~��7�߾�"�k�5L��B"��Z,��?4�2�ji�a2��� c3P��3/���n����E�h�iug�[���xle _��]`�ʦH`�7�%�>���+��H��(K��A4��G�3N�>%������"�6НO�{ڬ� A�{5(~�Tn���`�jh$,!O��b<C��g�0�>O;0FщG��� ���?����.�3/m��N�ü	���صZ�K�N�`�h���L�ޚ���O��k<�ȉ ����^>�u�+6~���;'S]�Zm��<塁u�<���`��i&=cW� ��3ќ�.�C�':fg����ܓ��	������j Uu6���c�<�'��f]U7���n>~$G���u(�8eF�gK��T����
��r邘cG7�D&�?�Ns�ŧ�W�%�#�ȍ�:<�	[��!ȍf	��Ө=�弈b*�B��+�)F���ϝ��Uة���QC��B=�'�����S��ǿ���}i�� 
G_k~�:p��ᓴ8�������;���E�m���i���S���Y�L�-����p)1�z}!���g,���1��i�l(���g>�tο0�S����_������~�ㆸ+�َ0���0��0��E�[��	lc�6��j���^���u�?��ZA_at��êP�B9��,�
o��iQb�F�Eۻh�v�Q���a���U;)P�&�2��^<Ģ�q뮸ȎY@����ZA�RF�y
C�@�s�(B3T�OΉa���\�C���= �A:wa/Dj?KJ���<ȥĽ��w3��m6'��Fo�.6:��틕dDHNb5���۾���4:�Ɋ��Kd���=ك7���^]E��m���lF�R��3B>�<�>�Qr�Ad��rɑᳺ1ЧS�N:��4Ny�Z��2*VUC�o��>ǿ/ťJs�]��Т���Sh��m��|�v"Mƿ_������<c �����7P�^?��m�y+:Y���k;���D�9$�)��7��8�"e�f!�O5��F�$/�-�^n�w+"�[�i�:��O���eIS5ˇ����ہ�_�T��A���HB��I�q���M���4������2\Bn\�6��c;��H'	�4~�`rB�������*e�-c���	u��8��[�A �6u���(m.��n�e_<��������p0)��&���~#��y�+�)��l�7M�7���d�]!D�W��|(΅
��r���3K_���%���̐�_��੎\y�x>я,���}�OWa�1'i�m��$+�;v�R~����
����L0}oI�2�oZN�Qsb�����r���ڟ~P�wT  Zl����h0Es�(�����f���v��"'Ф]�#�7I�kt�j�����c_�1���^�ַ�98�onNk�����e�KX�q�?��Dog|v��*��5��kh%axa�+���!��/��!U(!cH�H��)���J�r�k���7]�
!��q���͋�nǃX _BX�(��2�����ͫ�����f�Ux-ı�UI<�^�����8QJ��k�~���(Jb9pc��iQ�<Qf��,�V�����vM��&t� ��f4H��x}�Su׺����U����/8B�&bN�	z:�3�9�g"ע$v���nf3��i��!(��+l��W&����0u�m
Y�
�� ���������e��-�1܋�Eq}t�o�/�UEV�F�=�zU��ą�7��@�S����I�	eL<�^��1֨�R�;�H-ҞŮ�[�Q����N����6�	�ɾg��}���ժ\��u�����;	E'�'.��f�&�m�a�\Ay�`h~CK�|��S̜Y[;e�9�0���8�����H��|�����Lԕ<[*%^-�F�x����R�l^�#������@w�G�T����(�TM���F�A�7���mP5�(���2����⟂9�mH��n{j����'�XHE�7����Oz��]0w��Ⰱ��v�'\a#$�0k$���~Kb�4�W����X�Q��
[ٶ���AC�U�$�J���O�G8��>^��Z =�0�>��2���X,����,��v��F"�F�[`�4�p�ͤ���>��DH�Fx9�Y,�x�a��L�V�.,2Y+��Sk�J���(>gۏ�%��u�ui����E z��vs�U�����_�C
:����ZQ0�����&:������Jx;:�$��&�}�+ϴA�7�R|�x��F�S�����\��
u��bC����S��ge�jM$$�ay��D��sL�O�L����� �׋���yԴݏ�4a%G��E�"Q㢷����YI�=��^�cz�u-2�� ��_�x�\�"z�r��91e����]m.[��$�۵Nd�� m���5�٣q޽w�n&%m��Di_����������j�P�R9ݑ������-�0�FM������t�dϲ�����O�K!E|��&����:��3o��)ӒǸ��J[�<�ۜ�@��a�a�W{?�����i�2��?{���!��?�����cM�є]"��2����,�+%��a���������H�9䅺� �����d��}��`S��=S�9�HeZ������ɽ;%��ϻ��?#�p�23kTc�X�=�qhH ��SQ�$\za�4��(�܇S�Y�ޛ��-�l��	�c,��	';8;��%ct�ج,l	y����N�a_h�ɫ���e`�!�%y�� w�˝Fk�z����ژ�&uk�L � r�LD��`����?�2�3��H{t���u��\ A��U\����'(��=�yw����N:�����4ZT���^ݐ�~�&=�����6P���@A��ڧ���6�fjH����ڈ��L;��b��(�1(�֌��1������f�����&8����qЕ<ڧ1�������F���c��ȟ�C�����R�� ������X]��H�*J��t�������Hi0nٓ�}!�4Lܗ@��t�i�;��Д3�GŮ�YA�o���<4��
~}�ȁ���D��BcT�p�%Z�L5�5�Z���L���SX��Z�[�r9}�$)�ٿ���j��8�"��m����l����DU3Y�����GG����(�a�"J�8��L��\�)gl_��`Gh�EՒ��t����T���2�)c.r�����\!� �a�w��O����w�b�';�<}�n�[>��vw��ߛ8\���sS�K�!�2~<�V��w�Ư�n�MN����?�L��)��<��% 8ZT]L	6fܗ�X�V0
XV����� O���/k��ۓ��#�7G��������!�*�b��� ���<A/�z{����|G�Z�{�E�.�`�J���r=X���U㐚>�j
@"j��o���<֠�膍�]�p�Gf��ۨ�T�����d�#,�U0�O=� ����ƺ�s�������T1.z�J�[
	K#��[9�1 7�V�͑��v ��ɨ�t��o&@��?ě�����8�>�/9��^�����h�Qa������q�U��S�&�T�	Eg�DG��~��\#���!n;-��E�+���٫
��VK8�P�j�v��8�Q�#���:�>�*ٹ.���ާ�d�nq$�t�� >��������mR䚠�Yd�-/3[�?�������1����/��w4�f��������1N�T�9-�+KO���F�iR4Qq�c�S�'U\��F�ͤ>u�i�wO���h�������Ծ�j�ڙ�`s���Ɇ�Q���f�����?0O͇�Y/�,=Ns�� 9��-�����},`�u��@��&��e�Թ,�:��g������?n2�ދ��[%�:�[	�tg������)�����t~&`���|K�����%3��F�A�T*�!�cCJk�h(sR�R}��̃-��Rb���s�*A����>�h+��vt3#���lhɋ�yt#���4�KJ�sS>5��HsK`P�~�5Όz���n�ęR$��[����Gđ.
��O�� ���_݈1CAdg~�"j8��=����f�
ȴ�s��DFZ�)��C���L�e<=(k����rC� !�V�zhm%9���sԟVL�-��S>��}<���7%�<���K4��?osL���+n�Y; Ԉ%6��=[6!����� �zY�7�Mu=埯.ր5��,�$���{(f�q+�5�ֶG����
���k�A�?O�U�=-(j��x������l�I'uROD~"ƶ�=�sX¸�y�pI�nC���#��Y��H�"�Y��N1(��Y��U}OO\f���|Gj�E�Ώ=�mFbG�#�)/|��iOi���<�fxc�y7D�f�%+k��m�/���v�sx4���c�,B{�����b�Ӌ�3��\���ATXPP�����O������ܶ���&k�$�C-x?^����`�Q�&K��6٘�0;����.?$��<��ó���I���Y����&�����A�ՃZ˂Gh7l=%܋����Ud�M��]�݅c��K.����'=D$ivt�Ui1��|>)����st�Bk��Tx$�Wռ�a��l]�AÛKL�.M<�4����p�O�6��嵿슆%����!&�����v�x��M+��GT0�\�y�Qy+�G6��,<kjsoj�9�Q�����%��2.t|e��ZR���3�M�?:ݩ'��v6�w*� f5��=��+R���$(�n�� 	��7ĺ�I�#�-6��AT�xk�=�jaģ�ѳ���k�<�Vk��;4UO��z��:�s��/b�]�L4�)[�%f�F��X4д���o�o0�XH�,��V�H��
���W�B8��1c>w�m(�@i��Gl��zj����/=loNw�/e� ��
��.��)��Vv�CX��ϯ���h5�d����;:�Pu�?ZW�����LD���u	1�,�#"�l�X�pz�L�Wc�@+0v<�7x[���yg���;���SUh�-ǅ^��4��(yfp?�p�MdrZ�@��`�l�RK��+����"��p@cr#���<��O��:O��KC��3�DZ)��-�y�O�n��-] �CI�;ˠ��Β0�"VS�c ���[P��Z�p0���\���8�IXrk���ʹcE���B@�Jp��I,=��;ЗeM=���'��hX��KG�a�0bjC�3�w=��Z]��g�ڄ�bT�$ !���('Y ��T�a=�(+�3�%��A%���o,��FD�
P��!� 2��6ƣ�&C�-~�IM��V��is(./�A@4h��;�e���gt�mϣ���X;�k�kG.����r��8E����d¿�e�,�t2J�r��#:�����|[#�_֣����r�lv�f�B�Ҙv��Cv��'��~߷�� �>�6���u(���mI��y��e9j.�Q�0�ZUX��%OPRo���*�/f��]5<�w�Ѯ�T�pN��������t9N$�U�aI�-;�D6���
�H�o) � ���D�G����d�xRч^ͷ/���U�� �c~��E�W��i�X�J����t�P#KqȲ�5vx��p��Pc(}�/�=ҹ����@�X���̜vnfdF�ɖ�@7�R #�\�� ������E�T�� ��igr��3�4LU�W? y��d�È=U�4��c���AJ4+�����T�^+v�I��:������ >�r��;,ȼ��uO���ZG){���E�������1S{&WR�4�>��:eH(ߪ���V(!�O�;�%[UZ��x)'�-�y���+h��Fa̵w3��m��Ǥ�v�O�_���r�a��X�����V���>e�i���������a[��,��I��2]y3F�1��z�]��!H�C���{|�����Wt�<�ziz��"��bG��#��58%9����v=�Vԍ����KF��I�wF�Ne&A�E�%:�.M�� Z{�\<G>V�r@��]o0�p���E4v����Z0;�]�"j6 Ԝ�#� |*�-����[qA� ����x��M�_�}52��7�_ǚ�u�@��5!�� Z�A���u[����69a��K]�Y?p�����j�&���"�8�H��j��C�����Ej$c���.-!u��o/j��?cP���`?|%�!��3jߊ�R�� kqq�w�����dbƍj�|������=e����D�
������ _4��HZ������Z=���Q!�Iт���Y������\�5O�#� o��q�ǝ�E�����Q��F���y \+��Rݽ\�'Y#��V�d����Bc�7�S�{����:�{�[-�z���1ͪ���q�R�"Լ���]�Qt�ҵ6Ib~��� ��p x^"��'/⤰�}�?��/��t2I?�K[I9�E����n��ZXw]PO�#��S���RCw$����.Bd-m�M�kwbu>I�G#��n~u��Q�)�����º�g��,s�a�`����P�gk�8wG�o�:�'#}�\h�p{�L��Q�)Mc@_�I��T�A�+�i�����1�SX�����Gq���h?p�BM+8ޙ��;|p?SY�G�|�$��t�)�pjPaK���%Dh���k��I w�)Ed¡W����<0F!��c�7�A������R��
�쿖W����&VY���c	OIU�����ÛKߐP�c(��O�[��̇g�׍��M,H�	��E�����������%�������`K؞.�5���k��`�94���e�i0·���᫩��I(�ݭ����w�լ�'WwYݜrL ����G��f>Y�%��rR��<3Ӻ-.�Ti�o���Ή濒!R��DN��^{P别�k����}�coRk���}��Y�����b�/qF�1������.�I��$�=ba�c��ЦV��w%��=��g��-S_Vу�����A�j��GV0���J�	�4}�K:!֯62�(���r (=Dh�w�m_9f��;Y������+���H�o䀥wp'�uz�.�g�_s�Ł��˿�`d?�P�;SQ��q��kv��K[�k �}��Qy@Iom1 ��f	��s<�i��KSa:�����C
Ӷ��tJt�tlq�)f�U�J�tE7I.*ض�LN���oz�R���)u$�r�˷�M���6�;����B����$BX����徟��Ha>�lǵ�ԕKzB��	���9��Y��Ž~(���`������ ��93[��h Z�%d��{I���	G���7�~�@i(
����D�GZ���)���<���<*HA�����m���F����?Qg�]�}��m��T�!V!�_�5�L�������6Ҩ�8V������i�f��절���{�l�`8��mV���`6�{�	/T�������V��w#��y{�����"�5Z���D���?�̭�MQ��	R2ϕ?z���>x���RC��	"��;ɱ����o���q���ϙ)�ks:΢��$Qo��[��-�j��JP�y��/�_B5<���\�9]T����:{����;Y�;����z��}�ޚ&��6
��,b��j��=EJ��~��@�PA6��%�'�BH�(���K��6���kG� 30
�l��U<M~�GJNx���|9{��K�C��^��.]$�g(����k��!�y{�q�%~{��[��9�aa�δ���L>� �s�����KJ��z�e���W��MUɘ��n���wG6�t��x<��:����!"٢c�aj�2Y͸����a�;�n��3�I�
e�c����]#�ø��xd�����S�^�o׳
���?Q��wƟ۪u����.�	�۰�z�p#�V����Nq�T������r�!9�j��u�Ms�J���5�s����9�Nd&4.21H+�)]��<-{%�gx�����v�N)�ia;�X-N�(+���*��zK���kĤ3]��?���"J�d����v^#+������+V�DF'S��Lo2�+\ͅ�?�N�#�X��\B�TM1�J�t��*٧��=֒<1���v��D��	
�3׆k$$C)��}|�u�A�o04W�����f�P�Z��lYBɻH���p(8 C�ny�/��a�����"�ڕ�}�\�o��[~���S�@��	� �C�n�`���F]�x�,®�W��W||x�*W�%)v݅�2�E����I`�ׯ�/�(KS����^��׾���w�H�_���2XK��cxR�[1��d���0��|�����O��-jR(�2���>��'��f_.��P�)s��E���>_]���)J��=�p�j�-u�����Ƕ�Vۮ�=N�&�IW?����h�ܮRR�]u�h6RÈ������H�U��~V3ܳP{[��Z��4���E���V�$w�~�Z������U�l^�����Τ�8+�V�+��Zo�����dj���2P�uW�r���Ğ�E�S�"kmylR�'���-������@)-����4�O�|�whb�n��-�@D+�t���"�٨��V$���04�AH[��g)���vN�� �5v�S���L]�ZV�5�mh�O���k[43���>���^ى�l��CRP��2��>}vޭ�U��97��������s߃��G�	��F}���p[�v� n��Τ�/�`�r��Y<��SL�ɭdA��C�1�T��T#�%M��@�S�J+q�)��1�i�xQu�UEf�:K�b�a(��p�Hq���9���W�'P@4���y~��d�E���'��B�B-��Y���aƨdX	����,�a�#rB71��s�I��i�"���5&u��aӼ�x��I�ߚ��������sjj9���}0a��Ai��e=�V���n�i���ur��͂�aC-͑z/�e�*B�4��s�tw�iP���u^m �!�k���M�K�x
q@�RM� Ǩ&XjO'�xn��I�cu�bC�N��r9M\c���||�t���ҙǹr�#v��ë�o�J>�X�5]h�j���T"뤧�x0���W��~UE���{�Y�I}�.tՉg�O+U�L�#L��>ͫ��%��$��ѧV�_>�Kb�\���P��Jx��p�q��Ϥˮ�.������t��3��]#��ő����803��Y�zk��[� ᇕ`�o�rhlf1%55_�E�S~���}�Q�"a�����3�n��\qU�S؛.��_�T�q��CѠ����8��1�����F���w�h2��1�s��x�g<�i)z]fz�ABۙ���D� G%Mͅ����*�W�T�c�_�9�[iճS�ʪ>�)���6v�C��-���A$ޏ`gK��dg]?�M���d ��g���/��|X]E�>Y��XpMv��c��;6�a�FJ��h�t��Lp��}va�����Pߊj���
�&�c�0"���s�9��,ɘ�_И�������i�0�ׯb��:�l��-����&������[~�|���zhj�k�#J�&��, [5@ g�M#���vI�%˫��`��	��ӯ�W�o^R�5%E+2��#u�+���c������+���R)J�_��;�9n��HD��鰙	1&3u��5�2?�7עU�"P3~���n��u\\풿�/�����d+��*W,���$8p�A(e��*6���{�w9{x� �����5�w_κC%����[<���%F�F�:q»U=��Fjn�v�n�Q�c��J�.��Bl���:4U�N$l�c}�)����;��U'�z����F�5��\߹�%�:��1�ΰ.��҂YI��g���7��ջ�tm����qb�Pő��}����mgv?�B��#x�զvТ|��ǜ�	_�܃lBsܨ�d�W��(.��[�8��e�߫��<C9�VP�@�9+T��3�����j	�U�a��Zc[>=���'��ԝ���㏯�q�f�3��(I���{A��5��Fً��'A���c7-�0��6hH�F6qω�H^�%p̶V����f|U�P�� .�;r�K��CJp� ����1j���[��FK�B�Ty�ヘ&7׀�#��a������3�s/84�+���]n�f'��uo�8��i��ZA� �off5��j�4��Q���7�f�w!)H�7��Q��x�ߪ�z�F��YJؐ�]�5-pU;���(�п�7U;��ڄShJSL���w���h�G^���.?P؁4��ͶI��N��'m<)u�5�PF9���}����,�X��
N�m慎 BmJI5?`O��0~P������ٕ?�d]c:1�ݨ�e�� ��|[FeܛI��BG���P^3���H����%�l�$('.T�3���az
o؇�=a���g=>�c���)�FJp�S�nX)a�f�E�1��	x������H�7���?jo��&����RBG�b��m����H� �T�V=��B�9/1���l��o���'�&�.q��|�Pz}�L ���^(�J���6��3�$>(6R.Q��[F��cx�RCY��1�j�_��t.|�*C`��p*A]Q߀��|�%�t{$A��]��0��RJ����5��KGD����2�_��G��$6S@?S�e�m�sހ��W�ƏϛrD��H#�LUve^6�A	�kuf=�~4�yF�'�CP�2i�ywK]�(��Z�J�ty��`JKaT�<�)�!r�TH��g����<1>hj*d�&x%p�d��URb'Ï%���1���r��9�",��V���~�춄�z��X��������pt���Z�'��z�{Y��d� �.,<?�������]��g�b�����AJOߤ/}{�KnA>|���͜ ��ƫ.zާ]�w2U�[+}�޻(���E����Tˠ]�>���N�F';���x�N�+�))��b�q	>s��I2ѥ�������~;���>�g-V A��g��J.��i(���.���J��3dm`3�&:����p8n�����	�J`�m�.0�$l�en��8h�1��IO�}ӏ��؅4��P�Q�9���Y��KNn�X}s�vX��sXp:
�w/��
����Ѕ����*��ߎ�|Eq�2,'��*g#o����X�Ƙk�5-c��6�w
���ws�}{�=�{��ȿg���Nz0)":�ܧ7�-�qxjr��� �*�oi�$���#�%g<>�$a f6����l<�W	��p�c�k�wv�?�vu�K���6��WެOm[�EKA<'��t�a�'L�,ٟ��gW8	�t���hR��Αgl�_�t�ߕj�]3õ0abL"Ѽ[,O�K��� D*,Y#=�ΒB���;f��䒝M�h?�7&���2}�o����\9k����,���<9��II�j�Yo�.*bG�;Ä|�f�Hb"L��dS@&��K�#,��/Pm�����&q�#^��ʪN�>���ƌ[���`-�Z�o� �+N�9c�=��=����<����n���Rhc�X�K�ϒ�t�&�D��;�d��7���;C�xt��G,���&C��}k��L��ۆ��	��OØ��v@�H�WPG�)��@xW��a",�޸ب���䫆}8��P�&�-�v�+�^�NzD�g;	,4R���,���x��\�Z�3���X!u���왕��x���?"��pu��Q����w�Y��#G���j��nG W,r��x7.�
��:�.Zv�����De��j��u�ނ
��Qc�L��&��a����s�R'���.ÔNhw�O�+�9�S����W��6��"�Ox��b�0܌Jm���\�:���=�o}+�`��X�f���<�z�`���?WW׍Rw���l��������'����F�Lx�D�� ?�b-M�TD'<���-�?�c�)gA���H&�S�)tOfu��ԧ�B,���b>`ksx!���*�$?r��p�o=@�L��.��hHH*H ӥ#�Џ�J�%F���O�=f)�w�ɿSL�ʋ��.ɤ��A@A�V�^'�Tn�'S��5||�9�7?ޛ��Bܝ�3����h���A�YEl�+
B��*S�r��{{��t::�~T��\}|*�?ͯƤa2ay��Ivs��Z̿8A�9{
L����;j^(�+�� �B���e��.q	��񩔽N<n>8l l�Ir|*�-��2���f�gWF6b~ҩ�:i�#L�F&-4�Hks0r���@�V�@f[ǣ�kQ~�!��Q�&�j-�!�ʔp�8ڛ?2���'	���8W�^ܩ�l8�lpf�ʏ&�\�����e�k�Z�*ri��q9M�3��
q��K�p����p��pӎPf�!\�=����`�2�ciǲj�#HcM�;]��K��s�5�(u��y�|_w�2����,Ұa���F'�ǫ@�\.�
�����&[N�%'���sA���݂5ކ�;TJ:�H�v7�tZ�۠g|/��'Bb��,�܂�bY��#�SN���xF6�߉O':]��D�u[����:+q�{*r=������i He��u�wƝ:�W��vE�X�w�����+q����|]���j��k���g�[S������r������h-Z;����G��M�|�����$�Y�|�V��&T���*�C]����q�*z�O�˴Lw��9��v4T�;� �DSL�}t���!{F���y�;��r��:4JD| ����2"f�+jrH)�[>�F@Jlz��]��W�'>޴I������ }��Y������Z��q��x|�ji�s�:d@xx�QN�=���+�فD���Q���5�����ѝ��F�j&�(�q�c0-����Ҽ��<Ճ�;��*��ұ[���fF�!���@����=�`��2�D���x��P�b�8�'������hE�S�%$¨����E`�z;���5�\�`����n��:��F��޶��#~�z)����XQ>��_y�C���6)S��r*I�D�M�}��W uGr+�Z�,�.|c��ٛ�+����Qf�ZV�G<������k�k)�jWm��勖)\ s.w�(ovEZ8�]�YC��NR�J^�2`/ �r|��w�F�9BR�\�0)��B�~�C�R��)$}hsFү��G���]�?+�ȝF��4�GQ�D��۳~U�aǢ$e`%#6������cs�;R�9�<�H�_x֔�ȣ�y����� ����� }€6�,ZP��+�2jy�۩�A,{�������дzz����:�.�9wN��ҝI�ڕ��u	�7���R�X�􉔝����-�M�l����;����>LC��55������:���?�oU-^ҋ#�)wFWL5oc�2���i(d� �Sj��s�(�[�d��ӯ`���k�N`������@n�ʼ�YҤK3:�h��Z/��"!l�j����>f�X���ߖ'P[��	"B�돰E�3PW�z@Q�}�Eݡ��u{��|����%�eH�!�fU�n��M�B��u�+��|٭��`�=F�"TE�Q�s�R�,>������e:`Hl5R㑤B��%+�3�����a�%��l��Xl����7�Z��Gf����t��S��&,��#l����M,d�=�_��s���&cj6.G��4̅��8(F���~��V4�ء�y_U��fH������Fk��q�����867�g��V�	�`��ɲ�� �W<���ώ�o�0U(Svٟ3�|�bi�z��'�������+#�Nh�jMaR��0S�n�o��Q6Ӆo4���$
��� ����7�a_������)��g�����(O��������)��+�O8�[(td�n�``~��lA�:9�����%�����
�Q�\��Sx�z�F�+���/���
�,�g�/`�v������;&ݯ�D۫�q��*L��/+߆}����X@� ���M��5��֐�vа�9Q0���{�pc?!ѲW��(F�W9��ހ������z�=�42��V���LP��m����lY
"i�#&Hm���sTyJ1"R"7�����1�@�����~�_�HҭH�}�Ѓ=T,IQ