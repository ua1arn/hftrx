��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� ����־���1N<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR�� ����־���1N<��;��� B]�pE���	x]̃Dj#^Da����M� `tf��5�O����z����)�,�˛D��w���旴4�����:��@���b���$[L���Fj�A䵕O4\�p&!�ō�|'���@N1�w�0XL���t�ے����o��f?��n;�|-���g]��]�"+�7��K��l��fu�Z��"Rq����	��[B}9��O��<$e|����w'��1�:�Ω�[@�qR�� ����־���1N<��;���u��w)�SU��T�d�ǽ�*1�8�'�?�瑮��plJ�Й�m��8��r���t��U+�v��d���	u\��a(�m�Q� Q١Ӿ�$r�O��C��0�� �b�F���r�x!ڜg���p�+�8O �L#\6Į�E�=�&��D�[���(��h��CV�#3��?	M��y\XFs���RL�a)��N���m��~篟|�<�Pp�#R�S�y6�'
8�:r&@d�'1DK�5�#��ʐ�/�?�#}�{�
��R/�#3��j�f�ɨVu��7���	x]���~ВnK�k���p�C���|��X��0��F@�4%�
�V[���@��p��ʞC�ݢ�ep�O��"Hz��"��L�&Tj�P�6
� �AH��J���_a�M��RwM��;���`�(��h��$�~�MUs �~�q� \���T��U	�1�_u���V����*o��֢v��͒�&z��T�`�D�1�~�G(�����Pm�!=�y����h�}cg�I��O5 �Z��[H���1�<'"doB;sѱE�%2�}���3$�" ����f����m�!=�y����h�}m�#m��9�@���E�s-q��u���;��l)P�u��F"lܵ^�ZK�1Y6�k�8���҆�|n��q�ghY�_�X����J��Y���S>�m؆\�����d��.JKF�X��b��x
� �AH�O~=�̯�FZk ��U8�}�=n��vs!��~�MUs �̢���2���V��m[=��slc�/�<�M��}�������|���=�(��/A����;���m�!=�y����h�}M���_oH]���϶	����ę�u���;�'�� +��b)A�w�yJ�x;�������Np�,�n4_�����e68O�_��u��RL�a)P���6z�D�~篟|�sA�)#iZ&����8�:r&@P`��dpfVpb��#`^���w`q����u_��f0� ����-�l��c��=nB1�>�稅��m�!=�y����h�}�#�?�G7�Kq7a�Q`��̇����u���;���#x�d�f
�,�;�NO`�!%�qQ>B�~�e���rz�� )Te(�X��m�!=�y����h�}�G���Aj�}�aaï)ZE,�j�u���;�;N��;�Dnɴ7�x�r*�6��Ś�¢d���9��Q�Dd�(����6���e�V�-(�¦�����W�ү���u��w)�S��X3�����@��."=��	+;�'d$%MJ�Й�m�X�LGA��7�_���4�l��<u.�fa�Lm�>M�pʢ���dI״Ψ�w�Ua�[���,dԌJ�-Jdj�.n�
����k�8���҆�|n����:Vx�p*u��Uk�4�~���J�Й�m�T�#Ȃ׬��;�Ӏטw"iw4�q�M�4	�Y�����\�4�sƐ�hd	��Zk ��US����HU�6율��'�~�MUs ��y�Zk�Ž��=v �'	�?��["nq���z���J�鏈wƠ��ҿe���n �����SK���B c��(�U����	x]�<��O~���J�ޔ9����IOZ'����Oh56{�I"�c�q�CP�ba�(�N?0{l��wx0�<�·�
f��o V��	��y����/���RL�a)�G{�<�����G�/9@rk��O���@��<��7C��HM|C`r�3<0��:�.u��w)�S�3k:�(�-�~篟|���v���$2����E��j8�:r&@x7.ė)O:���?!Jf��`z$�X!{^d���J{")8�*I�����%̝��9=����RL�a)ѻtUWR�N	:.���n:�ƨ�Ob�N`�gը�d�7C��H.��T�c1����)zq�M�4=g���J��c�4��ic��S�O�4�B�!�6I	�Y�����\�4�sR���i1�����W)����VIW	I��?G�~�MUs +������\���T��U	�1�_u���*����	�����	����LO9� �Ŭ��2Dm�x]��.] �'9�����L.��6�H�.���2/�f��=V"N�^{")8�*I�ց��6 �����Y<�zd諒~����L.��6+Q)?^R7D�y�B.h�hC���(:�J�5`xt��R�m�!=�y����h�}�N�5�%����b�:q�7�<^}o?�M��;]A����@����P�����?��� �S��aY�@�Nq"Jc�l�!Hr�O��C��0��$�>��wަ����2�"�9����u���;�'�� +��v�ӫ�!NX�B���")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�;��i΀�cS���?@S:ӓ��|Q��&�N���.����'V��[��|D멼����@�Z����W�<����tТ���J/g���p��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"�4d�{!o�ѬL�1m��+Y#_W���Mz�8A�P�](���������f�ħƿ�9c�I�?g�f�Jm*)�m��+���qH�Ն��±�h�s�JFAa��Bzb;ym��+r��JʅY�y��
r�(����5�����x%~Y�1�:�Ω��
�/�rD���J7"�4d�{!o�ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l�����������fe�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`��'p�@�I�?g�f��m����bi�ī*�7�[��]�Xy8��;6aJVlO/	�Y���#U#��F��b��}'�U�4��X�Ặ��Ϊ���Jjz�^�R@Κ�2���ei!�`�(i3l0��F��j��#����j޽���Ǜ�����������i��Q�^�y�zL͊�q���Vǃ��������@���k��!�`�(i3�b9���j}8o{:��͹ ��1�Z���=�������Q�^�y�zL͊�q���}t��C��>�~I��M�H�ɇM��<
DN��b9����4�6�tھ[���:lw�0�=<MW�-}�	mp�EN��S�IÙ=�H%v@����fnQ�rV�ά���)"�,�>E����\�v���GAџV^�R@Κ�2'�̗������OtBl0��F��jT�����N��2�F�P��U��+�XhU��`��&�Q�^�y�zL͊�q��UG�s���Kǹ|���|u��R!�`�(i3JHn��z��r9�3�����$� �á��ٕ)����i3<�f�D���X���`	�"`��,���Q��K������E����F���8�TP��Vchw�D��y.���=��܄
)\Y���E����F���8�TP��Vchw�D��y.���eŞG�T(�E����F���8�TP:(�������f��[���p�ϵ�DEN�����M�*B�[zL͊�q��UG�s�����S2x�FRN�h��@���+�J��U<o^.K�}26U� �K%U���?�j�\�l�b��KQ�AF�E����F���8�TP�=5Y �������w�bk*�����y��|Y�
�}I�?d#De%�Ց$�'n�^0o���˟y��l�9>���ײ]�4<Ӿ^H��	�E����F}�=Ll�����&}0�@�͹ ��I�Q4p�/Cj���C�1��;�׊�:zL͊�q���\��;�,��yN4&�iq�VD�Lg�q��Dv;gJHn��z��r9�3���(��q�
�Bk�i�E?�xu�pW�Cy�w=�4e=��-�g)�X��Q�u������(�ʉ�I�,B�E?�xu�pW�Cy�w=�4e=��-�g)�X�:�G�
f����\{z.Ю;��!�`�(i3���+�J��U<o^.K�}�$;��션˪��/h�Б����!�`�(i3�E����F���8�TP��������ERF�G{؍��R��j�.(Wx*��|��pe���b�c��Et��q���U����?�!�`�(i3��|g�Y�'���Xw�E�i�m}6	��	Mk�rv�ј�"��Z鎬����A��:6])�/g\�H)��,vw+�ne.��xu	���S8����ٺ?��Ʃ��6��G"ڻ^!�g��U-�ee�@Rv����my$�N��o�/���;�%ؙ,{F�"�,�>E���TD��ό���.ӈ�=�$��zigzA=v)��(�
t�ژq���U��ꢤ�OgB�Y���c��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<������K�]2�y�Z鎬�������(����U6�bL��W��_�ړ8���/�����FZ^�u:��_x�����	Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/�I<��f��tN2s���(����5�%���(�-X�Ç�e���Hp�$-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/�7G��D�:`�'ࢯ�GB<[�(iN>�4�
�����Bdʨ,��偋:�Q	Q��|��Ӻ�(,��y�ӓ������ �V�ޒ֙f���_����}�\�����Ք�)�"JHn��z�c����,XL��=d��z��_#Ԡ�T��Ɓ��~�26��\�o�mW��y�ӓ��Dc4Ƥ S!f#���������l����O	%K��ͪM$յ[+8��"Ě��	s�_�5��ǈ�A0
��_�P[f���Ն gWVbT+��uL-���S8�,������9��
����	�|���/��@���#��M&s��'�PD������Y�L�FZ�1ǝ?nQO��B�f�8
��u��r��f���ՆnZ�va�?��Ԝ�G�ǈ�A0
����m���Yk���y��j��kj�����N��U���q��m"b��_��.V��(������}Dq�f�HN��R���מu���'�N�T~�m�ڨ�hծ���%>�rGO�D mWNHN��R���מu��� �H�0��
�5ߧE4��ʥ�nr]�b�N��?�{�XԲ���:'�>����߰r�n���D�߼
�d����ň�3Of'�����4�o�r�\Tȭ�3���r�<����M��_(����@҄���G��A"�U���w�c*��t+��I���XP��Ȗ�!�Rd=��¾ȼ�����Y�L�FZ�1ǝ?nQO��B�f�8
��u��r����َ�,�f�d��j�W'� h�ҩ���=�g[V��M*�/3o�U�r*A&-�Ri����l��M�r!�B/(�B���l1tSjv�!�`�(i3
ҭ�3���O���w�_f!�`�(i3��Ě�����}Dq�f��u��A�0�Ή*��a��2S����R�5ߧE4��	��x�(�6k�4d��!��Z!�;'�F&�MB˖�4,<��Ě���z&v��\�����3�}@��9�ڮWm�pi����Q$n�ti��|�@T��޹�{kb; ����ܕ����������a�"�Z�>)��]�B���[�.��|ȃ�$����T����i-}�����&;�8��������@|������]�^��� _�HN��R���ء�I����hڻ��:��L��O��݄�$��F�Ճ����\&�}u�i��|��
��(����{��ۮ�/���YЏs/�i���M4��S�$j���f����lNȲL���"��y�X�:�.�AY�@�W���� 2�AY��)��c�H(�亠-��fn�����I�#��Zb�JHn��z�c�����<�W�C%���6V���~�26��\�o�mW���'n�^0o���˟y��èV7�%M�����$j�@��+X>N�q�p�e6�_���|(�6k�4d�{j���d��,3y�@�VҒm�fF�5.]�����������0u�\k|aT��3G���(p��1Pw�������#p��H��R��Y��[�нx*�U	s����{`F�I6��M��^P�h$;���pM���ksdDH����'n�^0oq-���N>�4�
��,���Q��b�s6�d+��#	T�d����'3��	�;�j�"�[u��C@��AO}$|~�K��������� 2��L����ֱ�q������m�q�)Ў6dG��O����14�7'U�1�R�\<۳�<�G=}Id=��¾ȼ5�����}Y��	}�@�'�C%�-"�I5]l�����zQf�H����3bQ=�3�� �֤D�A��*ȑs��-�����y��j��kj�����N����"���jVѭ@;�jmT�#z&̴T	�et�f'%<7�lv���gWw��-����!�`�(i3�zk����\��;�,�Ra])n#���r������Aڬ&W�y��v���z��N���!�`�(i3�<�I��y�G��C�m�]6^�Y�ѓ,��|��H!�`�(i3)�{6�U���Ra])n#���r�����y��j��kj�����N�
\�n/S-��}Dq�f�HN��R��bP�63Z�tHN��R���O>�R�`t�td���5��Ě����E�i�m}6�E`���ʥ�nr]�b�N���pl�4ʀ���ߦ ����Rn�pPip<ɯ�nv��2������開k����6U٤!Q
���g��Vܙ��t�cُ�Ջ6�x�p�=����w`q��La��Y�E����m�s�*�MOL�ӯ.���w7G�����]\{���bq'���7ג��W!�͘�<�W�C%���6V���~�26��\�o�mW���'n�^0o<H�-��*{y���� �!�fLf��),��9��"!<���+�37y�����:���f���,�';:ZËF�3$����Vܙ��Lߝ-�Nr��VYW\-@��F~*7���&�_],)��v@˼�\�v��\aьIR=Z�˙}���.ᬵy��Nn"��%[��o@�?� Zh�R?�R��n�#ٷ�Ef��dט�w����j����r�C�M$�&d�X0�� ���3�ҺIÙ=�H��M����A�m�(����3�y�ܓr��G(h���i�K�g;�\��f9��NJ������@zLо$ԠI�*׿j�h�<�&d�X0���E����F�'n�^0o<5������U��֜��3��P=@��������$��Xo���~��1�51	�<����ry��cTx z�Jm]A�/����<.+6J!�5����`K��� �"�W�A�&hH\!�`�(i3�b9����lY1�ËF�3$����Vܙ��|�CY�oO���^��t���9j.�l>'�o��&L���W=D��'n�^0o`�U+�PA�5����`K~����G귈nIg�R���]6���b9���P9b���dט�w�����{�������}>p~z�r,J����!_�IÙ=�HB�q;�~ =����V��g��cH�wA�?��6a/�j�m��\�vňu�,�s�p�m~|��`.t��J��|�����IW�A�&hH\l0��F��j�q	k���A�P4ǲ I�g�R����z'/)�� 0�s]7�r޸��zL͊�q��o����6J��z�h��4�*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P�|h{�T��`�)�	�%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��Vx�%L��W��_�ړ8���/�C=2崝��b�7���U��+�Xa�H(�˕�%LH�N3���XP���f�Nd+l�Yҽ֗��D)�q]�i��E��T�
���A.o�G�m�?[���S��IÙ=�H��H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	���P4ǲ ��V �-�{q�����/��+l0��F��j#w���	(���B��j�Q��9�V�ݦ\�t!�ǿyXAm�� ��<��]��i�"�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\蟖�S� ?�0��E|�,°������R�wX���dט�w����j����r2��������������JHn��z�>�ack���A�;�֋`N(��/��<`�.M�� ��˽��r� B^�.�ߘ�)�I0M�/�s���'n�^0oPpkiq�o�H�MPq6.��[�#m}�
�?�A$�ʁд����-VL���+�J��Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?�A$�ʁнv1a{J�-���Ƚ�0Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�ϴ����-VL���+�J��Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�Ͻv1a{J�-���Ƚ�0Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�Ͻv1a{J��8�P��Άg��dT�W/S��8(�E���Kt���pm��)|#9���b!��u�ϟ��7�4�-�`~ ��#֫��/�*ܑe�W����n�4�{lGD�V�Bf�Nd+l�Yҽ֗�6��H��q���N�t�3���_���&#ݟB�E`^n�&�
_�n�@/%{�;����f�kN�ı*�7`����\Z��K��i3�|)sՀ�/V��������A@"�,�>E��k�:A�	S�r��AR1<]Q�I����踫g(�r�N�ǁ�f�TB��vC8U�@����gG���:���U?�G%ZQl蝌b�Bϱ��ᵉ3��鑘2����.0��jOT���hLP��2�q�7s�9���o��S8�/ #O�)�����}>p~z�r,�L;Л��|#9���b!��uፂ�6J�Ko��E�`JcU#֫��/�*ܑe�W����n�4�{lGD�V�Bh�5,Wlr�r%)cAh�߆��y�����DzL�ł)w���)]���&5j�d�٣��c�A�L'�R�M`Si�c�n�R�HM���#ga(􆿳�ټ*w2�56�
�CӞD�+5�4��c�%��)� BM���1�
�]�!��	Ǹ�y85��O�\�l$�L�溥����v�8:ۛ@W:���#���F]����.Zx�.����#���Ʒ��t���(�犽{Tɀ�$����nQ�rVt.�N���G��{�ݤ!�8���/�I����"�]�N��&�|���|��] 1�0µ�]�!����w�Հ�����DzL��T�B�X
��չ�Ad��d�٣��4�5_�o0b!��u�)���A7��M�����d�٣��c�A�L'�O�({���p~z�r,���^���2������}(Q6D����d�a�4$�b!��u��V����Pјq���U��@����gG������0w��z䮃��ġC���}�
�?�`)[�-hnqo)}>�	�ғ�vq���q�41&q^�`
�c��><�$2��Я�R�wX��}�
�?�`)[�-hnhG�W�ғ�vq���q�41&q^�`
�c��><�$��;mQ��8���/����,D��ǉã1Xɟw��D�A(g
�]�*��q�41&q^�`
�c��><�$2��Я�R�wX�ո@����gG�DI߃���iA'R�	�_��<��E����FZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕ #EO���h{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Be�)\���!�`�(i3�[�l\�`�|��K�z��@d��ץr�&U������G|M�Y�Q��*7b!��u��N�|�c�$�t�!�`�(i3���+�J��Y�{'%s�[�&B�踫g(�r�x�y�Zgl�k�������NI�:7�N�5�%]���a(􆿳���2����.)}���/�;���_!�`�(i3!�`�(i3�􇃬Tk�H@H�֦g�㎏qló��@d��ץr�&U������G|M��=����)}���/��C�x!�H�Z���,�!�`�(i3�U,�(�)8Q�y�� Y{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Be���`F��~!�`�(i37s�9���o��S8����ٺ?�n���㬺ƃ
ᾆ�x�T�\ ��i3�|)sՀ�Oi9L�:�k]m��y�1O�r^�!�`�(i3xZ��j�
�����1��;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J�O+T-rcs�"�,�>E���]�!��	Ǹ�y85��n���F�r�f�t���ӯIJ ��`y�����g�,P�n�R<���Յ!��4�c_����+#��.X���*"v%)��Qcm hP"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y����@����gG�DI߃���iA'R�	��.���E����F�R<���Յ!��4�{lGD�V�BnQ�rV��q�t7i3�|)sՀ�Oi9L�:�k]m��F���d H��(әxZ��j�
�����1��;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J���ǔ���'�P$��<�7��V�����T�=�;^�6#9���k��$a(􆿳��Y��$�	b!��u��Ɔ �����O�����PX�÷�������;^�6#9����!@�+ufw5~�.�.ᬵy�����3��
3h}Nw���85Zt�����V?�ƇBHx\�'���Xw s4S�'�i��`�z������ִG�ĵ�I7��-5��6��	���`y����@����gGI��l��i�g���:�a��Y�{'%s�[�&B�踫g(�r��C�M$�#ã�fޅ������ϲ�CyW�f�tR�wX�Ղ�hF���H#
ZM��L~΄gO�3����?��ҹ���+F�+�V��+�_��<��d�٣���������ݹ�0���f�Nd+l��p��;z���>)0'6���;8=�g��U-�e���b P�։-�.l?���݇�T%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7���d�uY�ة�;mQ��8���/����,D�I���A���]�^�kvo�Apw�I�N�_V�ܔp�l
d�R�.��On: +*��YN�ǁ�f�T���j����^��E���!��=T,��1�~�� �(׸���-��i��+b!��u፞�f
t斃����u_7s�9���on�-�6��
�jW��D���M���R'),��`��wu���뿼��8��''6���;8=�g��U-�e���b P�~?�b�e�2����t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z�����8��''6���;8=�g��U-�e,%�0g����A�YHm��G�m����E����F�i�_:�ܷ��	N^�U{xN��i>w��˪?�-�l~�U�n��(���(w�.#�U�EOEe�1<�6�n����=��H�Gc���=B<�O}����~�k�Q�)�v���|ۈ�٥��m��_t��:ʰ���w`qԴ�~`����vQ� ��}�
�?��,��	r�:M�'$�*��BL�Jx��e�2l��4��a��se�ξ���I��RhF���k��76�C=2崝���^�9�8pQ�J��7��!�`�(i3�Q�^�y�����9�!�`�(i3!�`�(i3!�`�(i3���Z1`�N�ǁ�f�T��	��S��H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	���P4ǲ �p�o*G��&1����L��h���vv���"	��� 2�I�Û[����N���gx$�O�Җ*���X�w�)?����t}�ݓ�ZeUM�ٝ�z*N�I�l�u������P4ǲ �p�o*����/�Z�k�ʆ-���t�]¥S��� 2�I�Û[����N���gx$�O�Җ*]��z�o̈�^d\�f�� l�o�bw��H(�T�O��{Tɀ�$����nQ�rV",�Ű�
iEE�G�p�o*��NB�D�u�y����R�`7�K����'3pk~��r�<Uee�N�����a"��-K8��C��Jqõ�偋:�Q	Q��|��]1B�]�b�C�r�X��À��#�P7��ŧ �GR��shbvk~�#xǩ"�4s2nQ�rV",�Ű��dט�w��^���֮�v�@[�JJ1��P�M��Ln��S�WY_���P[!�`�(i3!�`�(i3!�`�(i3"�,�>E��C.W26K�~�a�o�yai�7]����'�C}���� oI��RhF��r��,����g�,P�nv�@[�JJ혮��רc_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�9)e�AjL�E��w*�t%��zxa(􆿳��?ƾ�s��	��6��	����}M�l8�	
ږ�|����=%+]Bo�A;h�F��O�i���AԢ�a\�W__XOhGp�&���A�]I�3Ԩg��U-�e���b PbL}b����*���G��4���r�W+`�x�of'%Th�� �GR��shbvk~�#xǩ"�4s2nQ�rV�}!�@�?0����s�Y�{'%s�O��W��W���}���i�����dq�8���/����RY��Ɛ�<["��+�O�JT��8D��V�6IWJE�\��[�B�L�溥����v�8:��|`��'J�	�LÆ��E� )�&�VR5�����b�Bϱ�r��������]�Y����f�՜�T�\ ��y�.�`L�.@E~J��g��$���M�;�E,;��0����GI$��ǂcY�~�s<��MR*����%���$������ظ@	,���:�<�L�E��w*e�΢���v��J2N��c_����+#��.X���*"v%)��Qcm hƐ�<["��+�O�/�#��P�h}Nw����x�/�c�ۡ���Z� ��(HU�î�D�p�&���A�2��:�k���`�z��Y��),�B۸��L� s�j8&��f;�P�=��X��/D$�"��! Y�]�7Syv�J�Բ�������@d��שI4��欱���j���-+��B�G}ϼ 8���hy�`�w��v1a{J��ٱc����Ɛ�<["���܁�_�0�ΩyO^~��M����A�m�([}�@��L�7�b�����x�/�c�ۡ��F</h,魰d�/�p�&���A�&�ʜ��q?H^��2踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��<�ao����O����Ft��7G��L�E��w*e�΢���v�2��:�k���`�z��Y��),�B۸��L� s�j8&��f;�P䒡�3����me":l�n Y�]�7Syv�J�Բ�������@d��שI4��欱���j���-+��B�G}ϼ 8����n�Jt�g�v1a{J�=���c�(~Ɛ�<["���܁�_�0�ΩyO^~��M����A�m�([}�@��L}�
�?�^)�G�B�+�WdM4@��͒r��ǩb�W�[r��-�W.���g/��ξ���I��RhF���k��76�I����"��)׺������Y�U���i���@)�l��0�L�E��w*e�΢���v��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�zk���������XIb!�`�(i3GYs��$;���$���M�;�E,jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ�)׺������Y�U��3Y��P4���U�L�E��w*e�p�������
��M����A�m�([}�@��L}�
�?�u����p��8��V\⯜�'�,LFb�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/�Ӝ�z@����U��@at3Y��P4�\�7.��v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�ʥ��G�M��K��'�,LFU�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�zk�����>�P,љI� ���۫�d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�
�CӞD��=2���H��̣������G���]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/�Ӝ�z@����U��@atA�ᴽ��d�1�~�Z鎬�������j}�c��`�z��Y��),�B۸��L� s�j8�-D���(���!G�{s��?������H�^M'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��K���B�V�C��k��38�h�3&�N�qB���'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��K���B�V�C��k��38�h�3&�u�p���n�]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/��)}���/����ly�P�r��n�Ŀhw�)��Ov�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D\X��!��x�D�Re��BE�tU�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�t�,�NL}�="��x8I�3L�*}F�GYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8��h��)ew���m���BE�t Y�]�7Syv�J�Բ������sl����?r�<Uee�N�����H�OM��`�@����gGdR��Ƈ�r��F�f�J�v���+p���X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G3�+��m\n�v�ĺ�(���!G�{��yn_Fu�Ɛ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOU����q�f@&��f;�P�=��X��/�ب����b�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/��.������FD>�v��Pn<����X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G}ϼ 8���hy�`�w��v1a{J���MB��)p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u��@��A���k]m���r��y��L�E��w*e�p�������
��M����A�m�([}�@��L�@����gGG5������{��U����d�٣��c�A�L'G~��6�7;-;*�7��;mQ��8���/����,D�;����;�;��O�"���Q]� _�rs�i��@�N3,(�;^�6#9���k��$a(􆿳���2����.�N��+�j����tL������	�Z鎬�������(����S� ?�0��E|�,°������R�wX��}�
�?����Н���A�Y��|w�j<�lb�rs�i��@�N3,(�;^�6#9���k��$a(􆿳�P<t8��3����開�E��ч¼xE���8��w���ȟ���8�M�$�愉V�Sup�xg쬉� }���n4s1��7�癆cg3bQ=�3�� �֤D�A�f�8
�������&S��e	�/a��@�f���I4��欱���j����XN(�U�]���=�w�Ηե>���Q=z����9�r�)۬
�,#�����K1P��8?W!t��_A�;�֋`N���}J�|���|���j�)6)-
�5ߧE4��?�{�XԪ��]^)��\�׎w�-��8n$DI��'����0/ܤ�(g��V���[b�I���\�v�n��l����:%��Z��4��.�w}?�(��y(���B������P�I��RhF��K�X:��3����s�c�����gv,��u(q��Ϝ��*@&&r��]������4���8���i�_(����@҄���G��b�i0[����8|o����q,� L���,�F�?��jO���a�N����+���LQ�{p�uR�R�W�u)hZae;s9=3
���k��7)#c��Y�7#�xIQK*QYc����it	�T$x�����}�	76�&�� Ӗ�tJ��K�]���!E'�"�F�+��^�6,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����n�I��'����0/�e��9�S���ތ�1��\�v�n��l����:%��Z����}�%��@��I����"���_�Ps޴�ik]�7A��(�n��rs�i�� ��*b�+W���F�^�Y�7#�xI��;mQ��8���/�C=2崝�Q�gL#A=�����ׄ� a
��Vx^��\�v��|z���m��P���ݪ��*h���'�a+��tI�F�;���N%�:+W�5����`K��0)]��w�b^X�P�NI����l>o��|��>�*�).zVW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�pl� �PP��ƿ�c �B�dH�7DR�i�Ρ��˧T������X�p0�&�����Q�a5���nXZjwi�U���Mչ�����Y��n�Z(Ρ����u�PBxN��X*d��Uf�Y9��_QzMy㥁�hK�'�njVfV)~�`V%'�\�*�c�E#
D�@���b~��Z��=N��!�`�(i3�d�٣��c�A�L'J����l�!�+���LQ���"X��[��Q[R�7�n~�x��<�,���E�!�`�(i3�n`5�fK�\w��0]b!��u��չ���1|���Y�ǒ��Q]� _ό���.Ӹ@����gGWm?"<��_�S�
utY�{'%s��.|Z���I7��-5��6��	���`y����@����gG�[bGf�_�S�
utY�{'%s���'����C�`�/�t�KV*�3?�|��T�5�d�,WT	W $V��8���/�I����"�nx��hѧ�F��6��U,�(�)8���0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ��i3�|)sՀnx��hѧ���Nz�
���U,�(�)8���0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ��i3�|)sՀg�j*8a�.F��6��U,�(�)8���0y�	��sC��#���FӪ�c�g<�g��U-�e,%�0g���p+�@�����NۥUn����n{�_�\[$Q��
�̞��>�nQ�rV�}!�@�?0a(􆿳���2����.�t��������˃�Iy��Fp����f���,(���B�����(�犽{Tɀ��k�V\���"X��[��Q[R�7kѶ���� �oi���:FI�������b�Bϱ���w�K���1`��vߜ�*�l8�b(������#oM|#9���b!��u�],��%s��O©K���AԢ�a\��F�dHB�Fvͧ"�f���-A�¤�x.�Knq�z���a�R�wX��}�
�?������3�K�?\B�]q��T�ٮ|�,
���1��e0����yN��7��aq���E���ss�T�\ ��)�g.�F�_�u��Y'G-+;X����Jn,���`ό���.�}�
�?�ʬw�S��зq8�Ј'���Xw���,DH�v������g0TF�'�]�!����w�Հ㸮�U�M��	[�/��87s�9���o��S8�l7�EL��>0�1ۍ�h �=���"X��[�d�a�4$�b!��u�V@���gx2�n`5�fK�\w��0]b!��u��4�	��`��@��⋌�U2ރ�8���/�����s�c�����gv�h�ц� )�\�~xy�Bp��!�ʆ�In��tw�?�b�>޼�\�v�	�+�&I(&�L����6�{�Pe�E"���m�PU}������[��p#ِ.��҆�3�>0�1ۍ�h �=��h��a,JD�_�k�W�A�&hH\{UY�Z�[2�h �=�)�����g�P�e�97�i��'���L�溥����v�8:hJ�tV�nQ�rV� �L_K�*��M���R��ӟ-��NiघM�.�� �i�aYB��#���Fν��E���w�w:��y��j��k[:�ۤ�U2̥�0�L�p~z�r,���Y���hvl��9�h �=��l�I�SCp~z�r,o �#^{���y����b�Ա,��H(�T�O��{Tɀ�$����J�	�LÆ�c�9ʼ��$�G�nJ `G�p�P���� ����F��O�8�c{}�C���B��	��u8-�_��C`N�r7�r��#[��Y���0�ȷS�J���4�����\�v�n��l���m�-H�h�U�p�ջ�D�T�'��k$Y��C�9I��@��F��6�!�`�(i3y��Fp����f���,(���B��\���V#��p~z�r,�b��r�
R�wX��}�
�?�oj�+p�K�J�iN�S!�`�(i3�E����FAԢ�a\��F�dH��|c_�m��ġ��,�z���a�R�wX��}�
�?�Qw�$��Z��/�dW%�!+���E����FWS���
��ʅ�-`JX-�ܶ�0l�x����b�'Be��
������n`5�fK�\w��0]b!��u�v�A�
^^3�V�C��k�HvL)���	���hF�]�!����w�Հ�JX-�ܶ�0l�x����b�'Be��
�������+NonR[�q���U��@����gGP���Ʃ8/Tu�����_&����ʺ�;[��]�!��	Ǹ�y85�A�'5�i��|�����I�HM���#ga(􆿳���2����.\�#$�ÙAWfי�b��}!D̅����<!GO#зq8�Ј'���Xw�j�7��[|��;�ċ�lʥԆ�V��,ۦ�T�\ ��i3�|)sՀ�}l�����@~H��k]m��n�_��-����Q]� _�rs�i��~�g�t�qN�c�B���)%O�lg�;S"��<[$��`y����@����gGP���Ʃ8/Tu���Ŝ��%ٿ�j;�Jw�зq8�Ј'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ�}l�����@~H�k����`T�]b �!�`�(i37s�9���o×��̙�F�9 }�m�f�Nd+l�Yҽ֗��i�ܰAb!��u�v�A�
^^3�V�C��k�&�c���d��b�pAзq8�Ј'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUZ��| �Ɛ5�e`��9����dz����NR�p�'q�-��nEg�N>Z�k���@��b�Bϱ���w�K���1`��vߜ�*�l8�b(������l__�I����J�����g���R�wX��}�
�?�u����p�����+X��FJ���--f�`���$"�,�>E���]�!����w�Հ�b02�O�0�5G,��Gc#�T�Ed!�`�(i3��Q]� _�rs�i�M�����geE�vx���ƚP�& 5f��e�T�\ ��i3�|)sՀ�)׺����\� C&����q��Z���2%�ɛ'�F7�Gh`��@�����0y�	�l�f<Rqا �GR��shbvk~�#x ��M��.ᬵy�����L7�oa(􆿳���2����.+w�7�@�Af8�ٕ��(�W�!Ċ&���I�JZ���+�J���q���U��@����gG���U�\ʭB��2�k1�h�H��*�I�JZ!�`�(i3�d�٣��c�A�L'��$;-,�J�d�@q�2������}°������R�wX��}�
�?�Z�,��#�2
��e�������m[�LEE�S�_�S�
ut�q���U��@����gG��y��O���{�6�*F=ॵ��@xзq8�Ј'���Xw�j�7������1H}�ɐ��/��HM���#ga(􆿳�)�~��^�~�9�>��#�DZN7�{��|� �6+^=N%����Q�K�5OoL!���}/
;$�Z��"���t})�}�
�?�u����p�����+X��FJ���-��{�"�,�>E���]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/��+w�7�@�Af8�ٕ��(�W�5���^�.O¨�����+�J��Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D3�.%�P;˥�'ܤ",����^�� �YW;C��K�ŶT���d�٣����Qq�M��H�_�ЩI4��欱���j���~(k��V�Ρݾ� Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܝ�v�02+�j�V�-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcep�y�G/Կ�]�؈9ϒ<�3$d�I�v��]huP��/��~�_Y-�<���������dC�5g����w��N�KW����rS���,�[p�M����_	�#-s����J�~AW#��WC�ڃ�P ��*����	�� ����\�'7>�W��	2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�% �t=���GR�D^;d9ךp�+�n�)D�ʵ�b��6���6�� gWVbT+踫g(�r�N�ǁ�f�TpD��ZOU;��|B����ɠ�o���3�Z��(����5���ռ�j����)w�n��ukh��=��X��ϸ��#|S������3[�u8�b�ӝ5�T�w�%b��Gv����Y���a\Y����+���LQ�Ih uq�?� Zh�R?�R��n�
q8�N��ݚ�Н�w¹��<d�Ji�];���w¹��<d�,��L����+�t2�0�趦����'���o���a5���>b�eIG�5�}�]���p.0��I�![�Do�9�:|ܻ�*t����$�¿DĢ�WZ���q����k��,�:�N�*�x-�E��%�~�X���陼��"���t��f�?ǉ�=�⒍~��i����C��Y#ѥh�k�`���wӨj]h�|jع�D�%r�=k�Hg��iqk�f�?ǉ�=�� ߌ�ˢ�{��W�#�r��8�Q�z���`
 ֢��-���V5VM�dC��6�g��|��yp�(���z��l �>���Mb&�}�s�~���_F�k-��苇��Fe#OOJd֯��
�	?�<��&I�������=�'}�\$I���ҙ����
�Z�S$��$!��8�ZLN�	���gotY�^���d���!im�ڏ�q�Vъ�D��F_Q���
����M����A�m�(��8y�Ɋ����Z��!�`�(i3��Ѓ�\4]���3�dC���L�m��+�Z����y�=��X�!�`�(i3�,\ަ�It��+g[�!�`�(i3����$G⃍�����u~xgA���������6%�a!�`�(i3�gCu(o?C!�`�(i3�{#/{�p�<om��$���J�!�`�(i3��'abW�5�}�]���rQ�4��+�]�U��y!�`�(i3�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��K�^����\_9ͫ��Q������(���^�,\ͨ܉p����O,8�ݚ�Н�3Lv	̅���X;p`�(�����!�`�(i3Gظ0����t�%�Z?��<�ry^�
�:qEp��:��Zg�Hn7�(�!�`�(i3[�л���7��+��΢t�3����6�i��!�`�(i3{k�h�+d�/Y�Z-u�}#�U��X#�v�%2��;b�-�2�V��	��y��_�V|��~֤�s"�Dw\����,=��&(I��Թ�Ty�M���f�Nd+l�Yҽ֗�E�����+T5�O�%E#P.�`��ai�}#�U���b�N��z�+�ϸ�i>hw���k�:5A��pw�R���y�7Q{��̯�,=��&(�鑶��i�mJ�0�6�I��)���W�w��fD�v�H<��cBM�e�xڕ�!ݲ��_O�M3���� ��'�m�>�.ᬵy��&.=��;��|B���r����ϟ��7�4̇���>ZW�/�#+*f�L�t��n!�w(�y?w�R���y��0�J����hЗ
H�����2��E�.�g3Z�Ǵݵ��z�q�hW�k�Z]R�2�v{7!I���6�{�Pe�E"��*X��[��7%^G3�ai��x�����<���4���8ݭ�~r}�m�>�.ᬵy����*e@�_;��|B���r������hb���-�����j���t�T��?E-h��`f���s��6}���iI9�o«IX0F�M��hb���-�����j�ݚ�Н��r$ɓǃl[�Ƶ�1tSjv�V�Ո��+5�4��c�%��)� �#�K4dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�B� �b��!�`�(i3y�}�6f&rG��Hb� h�ҩ�V�Ո��+5�4��c�%��)� �#�K4�+�ϸ�i���U��[��c����l�}0�����U��[��c���@��w?�g��U-�e��:̘Ezł)w����ʮ��?G�+5�4��c��W������&�K�VF!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f���ܐ�}ī��K��M��lak���\�	�Z��.�g3Zv���� &�\JG8:B1+D?���2��E� �k�3��6J�Ko�.�h��>y�c)�h�<om���K���̂���Z��.�`��airV���qޤ⑗)�Ny������!t>rV���qޤ⑗)�Ny��?�����/��Ϛ+5�4��c��W�����+���*#nC��6�g��:�r���(�E�i�m}66j�"Hs��'o��4�Sf>���}nS�|Ts->m�9V��lak������t�T��?E-h��`f���sC>��Ӛ��S�J\7CZ�zk��Xl� u�<��DfQ���r$ɓǃl[�Ƶ�1tSjv�;�x'_|~�ܦ	&�P��ۥ�Y�mK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv�V�Ո��#�/=鴙ɔ9Q<ϯ��U�kSwgҠ�(�2j�y�`CrgҠ�(�28�Z5	Aݨg��U-�e��:̘Ezł)w������U+��_����E�ł)w������U+��_ �2���P�d�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��7���9iIk��/�\	"Ҹ�YlԘ=������	�+5�4��c �&A�5I��RhF��?�1�{� �k�3�?�����|2;$�J��7�OT�,h�5,Wlr�r%)cA�T%O^,v7�}�!��Tq��A��s'8��dA�IX0F�MV�ҁGG`5:��O.C�U��B��-���{�8�4���scX{�X!,xjzӝ���I(͂��-����!�`�(i3��6J�Ko��k��G<Y�dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�B� �b��!�`�(i3y�}�6f&r#o�]�ʄ����$[ʓ���U��[��c����l�}0�����U��[��c�����hZ?�JG��Hb� h�ҩ�V�Ո��΄gL;�uA|�d��Tq��A��sxGj@����:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;���z��O�3o����U�����0w�R���y>��yСQ=!�e����%.gW>�a�?�����U��)���Y;e�iK!���d.O.C�U��B��-���{�8lJ
۲������"sS<�0�zG�������&GV�Ո��+5�4��c��a��IN�ǁ�f�T��Ut>'L��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����x �͚lCv#�/=鴙""{��`j�#�/=鴙|A���a���1{&��� M?��y�!�`�(i3P���x�NSB���j%Ř�I4��欱���j�����Kk=�ذ!����#�Q���l�G�p�P�Jٯ�n
���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}Ę'w�4�5��ޙ�;ǋZ��E��3?�d���&�A��\x��;P����l�62�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�]DnQT3S=�t/�.A2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�@�Q�3ԯA?~va}�w�a
���˦���X��lM��m�w���i���Z���G�dE�h*M�jZ����1�:�Ω� C�`N��D���ÿ0�^��p=��X��ϸ��#|S������3[�u8��p�ϵ�DE�U����L��g�e�J�Pn\�}O�_�H8!�`�(i3������ET�zn�x'��݁.�q�0��E|�,�k�+9=�r'Z1p8 1���H-�`��E�ݦ\�t!�ǿyXAm�,���9^-���2��̪U��֜��3�kޮ��R�^Ƒ��f�?ǉ�=�]{��_G��JM�p�]3t�ݚ�Н���v��z�Nt����$�G@��@�D�_�k��V�E�-�9�ݚ�Н�EfVNNp"��R�ٔh8����Q��K�&�C�/�dy��7ht��}j���0�x��r6�>��/Zn!���ͅ�_�������� "5�]�/��@��.y���,��O̀�/�������� �mD��覭L��2��}���/�^��.@Kq�Ca����s���c]��H)��hy��)]W��7#OOJd֯��|��p8=�[Ǵ��p���@Z��
�	?�<�a�/!O�+�_0c ��X�\A����8�:�����zV���z%�/��Z>L�'��D(M&��7,������Z��<�6�Q=��C��iF63���ш|m�Q� �$^�.���Ԫݓ�,!�-DJ�@{a�g�G��4ee~1�u|m�f�<�6�Q=�q�ĉ�D>��2�0�+&���#XYKh�O��2��F�ΨM=갈���R'cf���8�>r&�N�����a"��-K8�T�\ ��;��|B���r����w��'�L�a�5@�i��g�)�I��#�r��8��ҥ�|HN��R��?�d���&�2��F�ΨMAͳ�bD�P-��ټsU6гd����Y)N�����K����F?�{_8�Y��=�}�Vݨ��}Dq�f��N��Q��ǺΕo�G�m�?���b�%ł�~�7p����nt=:�$r�t�}iV��	��yvѧ�_�.K`�J¹�0�
�pqPv�G�dE�h�	�t��������3bQ=�3�� �֤D�A�W�G��!?�d���&�x��7��0��jOT���b�S]O�lK��7s�9���o��S8����ٺ?������}>p~z�r,�L;Л��|#9���"(<K�'P�1r����:)�
�9�P��IY�]�!����M[��Ǣ}�
�?�G��-�HG(��J��� �a2��*G�� ��x���rs�i��9˹$m��U2��53��MN�-���8���/�dТ���S�d=��¾ȼDw\�����b�S]���З�^���H> �a�{°���v1a{J�_AA^_n���|ʡi��!�`�(i3!�`�(i3!�`�(i3V[B�5�mm�ڏ�q����v=NWv�A���U��)���Y;e�iK!���d.[�����:Fa�7�����~�L�>��',�$R�i�Yl-��<���xjzӝ���I(͂��-����!�`�(i3��j�4�<�..�4���J�c>�$�my$�N��o�/���;!�`�(i3G��-�HG(��J��� �a2��*G�q��<��K�my$�N��o�/���;
�:qEpk+Q�h'�Ȝx�5W ��̫(� h�ҩ��H����o�γ�ha��o���H�RtV�^Dw\�����b�S]O�lK��C&��b�:)�
�9f�!�Wm���m�q�/���e���WƎ@��w?�g��U-�e�F}�.S+t�Y{�<����
�9�v!�`�(i3�T�T�y����O9�(UҔ����F��l_|�(��j�4�/�0���p15hQ�SQa�dz��q�+���xҩ��ga@MxW�iGw{z���"X��[A84Ы�"��m�q�/���e���W����^dE���b��Bg����;?�P�d����%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M��ŊPT��b��Bgj��i�s�)�{6�U������m��U1�� ���zg(LfÁ��/�0�I�k��q��־G3�ai��[��*"����G�������������q� N�}��������Q㬍�G�dE�hi��7u�`����k!�M�Z���	��51�X�c�rs�i�}�O��LTSG��ʎ��ߜ�2a\c0@Ɓ��"�C�ף��=�^݊��>��B�K��b�S]O�lK�������[$R�i�Yl-1�*��i��ċ�!1���~!�`�(i3!�`�(i3!�`�(i3!�`�(i3=��a���my$�N��o�/���;V�Ո��!�|_@��0]�9�x0zޚ+5�4��c���]W&m�ڨ�hծ��.J7h����}y�U�@�stU6%�DK��\��u�Y�KG�ξ���I��RhF����u�*��?�d���&��ݚ�Н��e�<Q����ON�C�'�@�E���N���U���H^�N���������$���sC���X)�{6�U��I��)���W�w��fD� 4� IkwqE1r-���#ȉ��%>�rG6j�"Hs��~��-s�*��8lx�~�����=,��G��z��/{j��06�!&>��q�+ �Ǵw�T:~�Y��"��5�O�%E#P��.J7h�4���>eC�r�&U������G|M��QVu'�e��0�U+�qbp@�!�`�(i3�ݚ�Н�&�z���@hӛ�/6��aW�/�#+*f�L�t��nWIi{4D+G��-�HG($R�i�Yl-%�z(�~�:)�
�9��3�����1{&��� ���jd�	�!�`�(i3!�`�(i3!�`�(i39�{�Jj3�8�`�`�6f�Nd+l�Yҽ֗������1xL��@�a��<	: � �&A�5I��RhF���k��76��wiV7Q�h�J?�߱}'��)I�y���j�4�/�0���p15hQ�SQa�dz��q�+���xҩ��ga@MxW�iGw{z���z�t����q���<�W�.�P�	��
�Q�}FwZNE�����A@�Q��ǺΕ}a�/�kj�>� {�}���my$�N��o�/���;���aR�!�`�(i3� 4� I��t���R���$���R��2�"���nH�W����6�~�5�O�%E#P!�`�(i3�mp"�o��^�+f�λ`,9�H�W�Q��ǺΕ}a�/�kjȍc�==�O��V��&�J��:����!�`�(i3&�z���@h�iqk�W�/�#+*f�L�t��n!�w(�y?
�:qEpV��	��yv�ʯʗ���>���}Dq�f��.�g3Z�)V��B�1j� lL��!�|_@��0�Wrx.�7ѝ�.J7h����}y�U�@�stU6%�DK��\��u�Y�KG�ξ���I��RhF��K�QU�?�d���&��ݚ�Н��e�<Q����ON�C�'�@�E���N���U���H^�N���������$���sC���X)�{6�U��I��)���W�w��fD� 4� IkwqE1r-���#ȉ��%>�rG6j�"Hs��~��-s�j� lL���C�߽�|휗��,�ǰ���9kn��CX0��W@^��}�Q�� 4��/��t]�<Lz+M�ᴰ`�V��rU�w�⽒��8�>r&���R�}vJ^�9���x��;��|B���r�����g�9��,Yb�;�
[�&~����w��FH0M�F�r�f�t�ŝ��X��MM
��,=?�d���&��ݚ�Н�N��	�Ȓ�@{2귑�'=��!��b&l�t-N�Ɔ �����Vd��0�| �艅�%>�rG6j�"Hs�ĖYS��������}Dq�f��g�9��,Y�����9C��K�J���֏^�M;�¬pX��D�P�E6�k��q��־�W+��W��G�dE�h���|f��ӡ`��R������s��ꬺ��1��:5A��pw�R���ykb>���p���㬡�xvrCw�R���y���,!�뱁�c
��X��u��V�H��;_��8W�w��fD���}l�g`���U��t�i��˦���X��lM�Ҡ�N�����?�d���&�C#/<���q�*���Nj�MC�%`zI\��!��6j�"Hs����]��.d`@i����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcזU!��%6��6!i8-0)��0�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���i;�Z����yQ�H���%�#�o����q,� L���s��$�Z;��|B���(��m�Q� <L��-�Mφ�q�©��ല���?�;��XC5,�����t�iZ]XF�hx��G��!�`�(i3��иܖ�:�>Xn6��M����|7J���U�ݚ�Н���v��z�Nt����$��U�좧���h �=�f�?ǉ�=����Kp&�@���k�֢F�7��Y�
�cc�V��ݚ�Н��כ��p�'��5��s,ݕ����׋�es��O!�`�(i3�d�uY��a��ZAδ�W����vcyj;��q,�zg��p���]c���H�p��@L�0�وݑ����1I^��+qѭ�+g[��y��j��k�lԇ�-{�-��i�m�T��!�`�(i3k/�z�xEQ!�`�(i3���*[UxG!�`�(i3�չ�Ad�!�`�(i3z�Gb��P�!�`�(i3�<��>��%@��4�䏄�J��9ŏ����V?���覭L��.J7h��r��H�:S�.?<����0�9�dt0j����i��NU�q�\E��0	ozqPD���K^�)
+[?M�y4����u_+�_0c �bYގEV֗�<�MP�>�n��-�U4��\w��˪?�-C
2��>�q;Rm�5�O�%E#P�F%�X�Ԝ�v�<�$��	��#4���Śi�׿j�h�<�H��q�/���˚����Z��!�`�(i3��t�f�2E�B�ӗ�z�NE'#�~N2��IET'=��!�̫z�����	HN��R��?�d���&�g������LksE`*@HN��R��?�d���&�zY]�埅؉��+�Ws��h�G��;_��8W�w��fDa ��^�0v�6���^�F��a�u��ݥv�1.�)����x���	R����>�R\�!s�A���_r�e~5�O�%E#P�>�:| �II���؄m��+��jTʱ�8F0_H����=1��\����L�,\ަ�It��+g[����=�-�o&l������g����=�tt"���O�����J��a�U"����N��Sx�M������p���,��2��������")d���ݚ�Н�Q١Ӿ�$������i��X;p`��ļަ��P'b�be`�t!�`�(i3ct�:��RE��]n��X&|a�#�I7��-5��5Z��=��]zŎd>&�&i�������kޮ��R�^Ƒ��f�?ǉ�=�B�6�N@���k��-��W����vcyj;��q,�zg��p����8��'@���k�� tZ�u���ߘ�)�Ij;��q,��z�_�Б����!�`�(i3�������a����"�$,\ͨ܉p����O,8�ݚ�Н�Gظ0�����@;w�$C,0�?��ʝ�hy��Q�#<4^�>N0Θ��ݚ�Н��ƿ�d�����&I���m�
��,!q�\E��0�����?Oǖqo�_����m6(\�]���f�?ǉ�=W����GS�*;q�j,���-�}s�Z�|�X[�m����!�`�(i3+�uB;y�L�6yd(�~��rͤ;��krk�ɍ���>Pҝ4��/��t]�<Lzg��<�=Lk��D5�|أͽgF"?�Q��ǺΕR'),��`�C,;�m�~�?�d���&�x��7��NmyM<�G�ۺ�Ub�!�V��u��i�_:�����k��$�8�B���ow_;O
�J��:����1�����j��G�m����t���[����<���/�sLXNAA�����}Dq�f�����,�ǰ����������^�)ߋ����-V��	��yG��Γf�-I�p��g�`ks�F���;_��8W�w��fDy�^ecK̅�8�:����	ڱr&�zbYގEV���{����/V��rU�w�⽒��8�>r&���nH�W��^�̷ؠJ��:����g������V���S����,vQQA�q�m�,�5�%]����8�B���ow_;O
�J��:����w�.Y�[�����V?�_.��45�$��cז�!�|_@��0,���1����,H/������,�ǰ���������{����/�_��.���9�Z�y�6nZ:ӄ��8�|����N!�֏^�M;�¬pX��D�P�E6�k��q��־�W+��W��r�+�����i�g��QZ���>�ĩk(�CQ��/5U���F�SRTpI��)���W�w��fD�g�9��,Y��(c$�,w�R���y���,!���f�|�H��4O��A�6!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc%�o�T�*9������ر0%W��2s�1��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcf����5�CX0��W@^H���%�#�o����q,� L���s��$�Z;��|Bq�D�7�P-7�vqq��R'cf���³5��*�7`����\Z��K��qb	��G��W+��W�ƻ�.=�+��T����oGo�Z�������/�)��ɖ��>��O/����Lt�iZ]XF�hx��G��!�`�(i3b�ӝ5�T�w�%b��G�
�Q!}-[�J�� m�Õz������\��������G��n�����������Zٲ�6׿j�h�<��k�+9=�#�-�p��8������aP��k�= ��j��`�3J�V����U����\��,&߰��U��f�?ǉ�=}Eo^��Ŏ>s��Y�&�������t���c,\ͨ܉p����O,8�ݚ�Н��$�`V1���n�|����Y�{'%std�jk�"hy�`�w��v1a{J�	ϙR~�D`�ю�[�T�tV�ǃ�(�s��0�;�l]�a(􆿳�+�'�hy�`�w��v1a{J�{���Ob�� ���t�=�v��*"3���'�C}ߦTd�n�g��U-�ew�K�H/�</Sn��'B�ɏ��]�!��	Ǹ�y85���J�%��[��m�Uƌ0Q_,�F�dH����y�����/��b��7<Rnnx��m��M��ٌ�RnQ���_A[��m�U��'�Ѱ���w�K�R he��as�C�G���-�p'�"�hPW���[fS����6s!�`�(i3���S�|J���^���e8�W{�
�s��wӨj]h���gX�L�m�;����ॐZ���*�7`����\Z��K���j�ONX\!�`�(i3l��A-���:��]]t|���|��m�
��,!��hy�NzK�}TR��b=�!�`�(i3�չ�Ad��vIn���9�Yt6j�"Hs�	��=[Y
�
�z7i�.�g3ZCy;"-����U(0�
�pqPv2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�ٻY84��s~�~�7T|2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���b�s�D�.�)����x���	R����>�R���mK�g+�Vr���J��:����b!��u���t�f�2E����u_7s�9���on�-�6��
�jW��D�: +*��YN�ǁ�f�T���j����g:M~�b1�Z���=��L;Л��|#9���Ă�m�DsQ�V�r[�}�=]X���1�:�Ω�յ�'�)xE���8�ب���H������%kR��������֢&@��&��k���t����~�.U�G���/��q�Z�n&f�Nd+l�Yҽ֗��ZE���n����������������i��X;p`��d�uY�ؤ��E���v:ι�Y+W���F�^�Y�7#�xIvє�&������0/�e��9�SW�Ty��5!�`�(i3���0/ܤ�(g��Vt����$�����p�><{ �=�%��ʒ�!fsZ�_�������� "5�]�/��@���Lt�2�t�&8�,������	�;�ݚ�Н�h�'f R!�`�(i3>N0Θ��ݚ�Н��ƿ�d���!�`�(i3M몴PBoT�ݚ�Н�?KYC'v�����#XEXj�.�nX�p��"��覭L��2��}�������K-�����*��$�q�ʋ2�ZwŃ��t]�<LzKj�`�|\{ف(�7�B
IQ�?X�,�7�%�a�A�m�(��X����_��s�֙7�}�!��ۆٗ��NJ`@���!��#�)&�-�y]/�qF�ŝ��X��MM
��,=?�d���&��ݚ�Н�H���7Ә,�۞��	�����p�?˻�M���foti�J"�T#��(�&HN��R��?�d���&�ۆٗ��NJ�F�}қ~Ĝ���,�ǰ����
k�=a�~~��z}�G��6j�"Hs��I�x�d�[�Ʃى�6����O���5�/���[�Ʃى��+�@t�L�FZ�1ǝ?nQO��B��N�����?�d���&���5�G
my�/�8yv���}J�|���|���/Q�������d���!i"(<K�'P��6]~T|�nX�p��"��4���#�`���m�jp=�>��o�
�v�ξ����l~�U�n��(���!�E��]1�Z���=��L;Л��|#9���O.C��������m����!(��'HY-��Yk"1/]���!E���VG%��v�/R�R�7h�,b0V�u�Q�ݚ�Н��������r�E�Y������i��tt"���O6/��������рӚx�f�?ǉ�=�]V�H7'�R�^Ƒ��!�`�(i3 tZ�u���ߘ�)�Ij;��q,!�`�(i3�z~~�Y_" �g8YwU��֜��3����d]���GF��a�1�Z���=�,���9^-�S�_�p���it	�T�=��?�AQ�0GȨ��_�\G�k�y'��af׍�Z���e����kn4@Q�/�!�`�(i3̇i�d�?�!�`�(i34�0 L?�p���@Z��hy��Q�#<4^�-����b=�!�`�(i3�չ�Ad�!�`�(i3z�Gb��P�!�`�(i3��TBd��pS�*;q�u��&�o��n<���AV2��O}�cD�����m�wӨj]h��
����ŗ&8�,��ĦsW�0��Ϝ��*@&+�_0c �X� �Ĭ1�<^��0�u"��D5�|أͽgF"?�Q��ǺΕR'),��`�C,;�m�~�?�d���&��ݚ�Н�ۆٗ��NJ`@���!���ƫ�P�A���8��''6���;8=D�P�E6�k��q��־�W+��W�.5o�fa��N����Qѕ&D�a�Y��m�'�¯ԙEI�s+��6�.|th1�$�g�ݚ�Н�w�R���ykb>���p׮Miz���;b�-�2�V��	��yG��Γf��Bp����ӛ�i��.}�	76�&�;��|B}2_R��'3x)'�V�*�?��O���2�"��H�ʱˡ�ۿ��j����H�V�7�}�!�����*�t��v+�/;$�������1�1F%јI$r�t�}iV��	��y�bB�.�����	7?�����,�ǰ�QCT�"�Ʃ�A���vA#&��Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�:1j�=�+���u&Z�=��O}��� 3[Hn��Xa�����`��O��m�]wew1"G�6L_i��Y8:0nQ�rV����X8(�K&'3����G��-^/s�B`@���Uc�`X�,4�?n�J�����W���h,3
V�R���S�sq��u�����|S����	��rc����	:�¿D�?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�{zY����b�8�dX�↨q�©����y,�m��M�5��=��X�t�iZ]XF�hx��G��n����������������i�����d]���GF��a�1�Z���=�,���9^-���M���R��ӟ-��ZWq�ߑ|!�`�(i3̔`N��?�R��n���Lr�VU����*
��c�<v���G?d��A ��+���LQ�f�?ǉ�=��h;e��w���U���І��%n3uZ�v|�E��n^���+qѭ�+g[���|��pe���b��˺�Q���f�?ǉ�=k/�z�xEQ�苇��Fe#OOJd֯�|�)՜�4-��r��gGr�����rk���6���
|j	FQ�)HVi�p"���#?�q�\E��0M7$����1Ʌ�Mi��������<�ry^�$���]׽��X;p`��D����m�c��o�;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��`�����J2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���L���Ŗ6$\K��p�>&�+���LQ�����_��j��N�֞q˩���.|�YtA[���Ŗ6$\K��&b���E�vL������ur]p�+#���&�x�.E�FY��+c��8���ݔf�zE�񪣘yg�U�։�������� h9�=�^�a�	�ӪЪ�S>f}f�Y\%wj�j2�%�}W���8�=�w�����5�O�%E#P��_Ѭ�Q�vC��Mi�ʷ��A�21�ri��WH�1�:�Ω��maC�S�s9ى�^�����L�,\ަ�It��+g[�A.e�@H��R�^Ƒ��-��IR*�fN�W�Ty��5!�`�(i3U����z~�B�wj$g?d��A ��+���LQ��(#��3��G�K$xE�p4rqG7�&�C�/?!���l�~�y��(<�Qp�P�N�I�Q4p�/�;ϔW�����1I^��+qѭ�+g[���hy�NzK�}TR��b=��y��j��k
e�3+{�i�m�T��!�`�(i3&��s���qFҠ0���g�ʈ�/�q�\E��0��W�tȇa�^��D�f�?ǉ�=D�wP�/�w,���^��5�u:/�ˇ��;_��8W�w��fD7~� ��Gs͟;)f���SS󵭆�ײ]�4���yٟ����_r�e~5�O�%E#P��Q*���j�va�>]�φ��<�6�@a� ��fFMqlgd=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^2W���R0�	�����e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;��l�'-�PM?��y�!�`�(i32W���R0(|v��t�a�^��D���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M|]η��q��_N�����,�ǰTm�v��G�jq��vĪm2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h߫G��*%\&%�=:���'��-�3��#?1�U���gFck
���&w��U,L���w
�kVr��)` ��d���!i���QB,�Ϙ�h��'܍|Cy�IX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н��lTN��IdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H����#� �,W��5��t�����F/G��Hb� h�ҩ��H�������
q<O�A'�u������O�g)�X���2�-��1tSjv�!�`�(i3�lTN��I���q�}���{BO���5�%]���a(􆿳����^��
�:qEp�;�P�t�5!�`�(i3�$���"�U��I�,B�E?�xu�(ݖ��Mb,@^;��u�u��r��!�`�(i3�du��m�_�3��+�uB;y�qT��#zɯ.�]ؔVG�g��U-�eU����z~��p�~/r����*�
�)g��ϒ��{BO���5�%]������[�w3�_�]!�`�(i3_!4rd A�_�3��+�uB;y�qT��#zɯ.�]ؔVG�g��U-�eU����z~��p�~/rP`��� �)g��ϒ��{BO���5�%]���%�gg�v���x��y�o�!�`�(i3�2��}��,3@97��jsrCm�k�U6�bL��W��_�ړ8���/���}Dq�f�՝� s�#���k$ !�`�(i3�;�%�R�����0�u8�a%�R�-�w���+_�mS8<�n�ݚ�Н�!�`�(i3�lTN��I��!���c�A�L'M�M˫ɒ}�+@2l2VQ+�3yK������v�h�Q����0�&�����ݚ�Н�
�:qEp'{w#/ B!�`�(i3q�\E��0��@Z���rs�i�}�O��LTSG��ʎX�����j�5�%]���"S�`�6�1�Z���=��n��I!�`�(i3$f��_Ub�F�S�1 �
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;���^�#�nQ�4�gX��>`���^9Z���;��|B7/#(��E+�g�BV����01e۩cS�e����k��$A�h��+Fen����9���(S˪�Z�w[����Vr��)` ��d���!i���QB,�<(U�}E������"?��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�?V��j�cF�l�q��my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�6��J��c��T	�����Va�ir�Yu�������&G!�`�(i3�lTN��I��!���c�A�L',� *�]�o/��@���J��6�d풪����R�^Ƒ�ӆ�v�9��HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ o�n�J-8$u�Ӵ-�aT��3G?�d���&��K"�d�Ҽe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�oA؈�'��(�.P�^����^2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�/��"p̶�X Hz��0|VO�⅘�φ��<�6�@a� ��fFMqlg��èVxjzӝ���I(͂��-����6�ZV	�	�F��6�E�g�������(ӈ���m�r�������8�28Y�^V߶�h��,��Aݖ��"��#���Ff���'�T�n��a�^�y��� �s��c��̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l��MmN}4��)j���;���N�B܍���� h�ҩδ'.�T���Bf���T�n��aο8w�B�Ra])n#���r����6�ZV	�	ҙ���˦G�K7͍��|��W&":�ݚ�Н����F��O��ݚ�Н����^g�6����GQ�kŕ��QH�RtV�^6�ZV	�	����GU�lP4����G�Ε>�E �Ra])n#���r����6�ZV	�	����G�^E4+у��b�Bϱ�nQ�rV��q�t7����ʻ)�	��-M<j��.#!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M�&O�a��B�5�S�H��ԻR�Z���#���2=��h��IX0F�MV�ҁGG%4vkz���յ[+8��r$ɓǃl[�Ƶ�1tSjv��Z T��F��6�E�g�������(ӈ���m�r�����Z T�֕�Nz�
��E�g�������(ӈ���m�r�����Z T�����GE�g�������(ӈ���m�r�����Z T�����G�J�c>�$�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l���oi���:�첗;|8,}'�%�y�ݚ�Н������3�K�?\B�]��*�·O��NۥUn�'��L�xt��s��kQ䖬n���S滑����ZLN�	���:����
�ݚ�Н�X19�-.|}���˃�I�xF�oͧ�ߜ�*�l8�b(��MdGN���!�`�(i3T9��JG��Bf�������3����#�=3!�`�(i31���~!�`�(i3�����3�a�E�Rq���my$�N��o�/���;!�`�(i3���F��O��ݚ�Н����F��O��ݚ�Н��)E�Y�ȣ�NۥUn�����D���u��r��;�jmT�#�����3��vI�o��v��ONH!�`�(i3T9��JG��NۥUn�J!�\���9mh��n`Ӝ�*�%!�`�(i3�����!�`�(i3�Z T�����G�^E4+у��b�Bϱ��L�溥����v�8:?�'��៑fI�[ ;N��L/����9>-WH�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�"�4����{�=0+�{�*&��q>�<�'���I����� ���JH����8����F)�~����H�V�n8�A�A�y���6���#¯��TG6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3�4br��n��>�my$�N��o�/���;�B�'��a�S���%��3|v��Eb�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^%Q�[�J��]�U��C�|J3J�W���b�0�;�jmT�#~��F�����������yN��7��aq����i��oZ O\������U�._�nQ�rV��q�t7�B� �b��!�`�(i3QV�=��̟�1��M���R��ӟ-���J��RQH�RtV�^!�`�(i3�4br�����zk2��/����*Q!�`�(i3�	��x��ݚ�Н��B�'��a����aGl���nF���<�W�.�P�	��
�Q�}!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�kv޶Gl�f��1.Xw�R���y>��yС�|ʫ��ď����~͏��{KH�"D'���I����� ���JH����8��#I�ND�s���H�V�n8�A�A�����aGl�n�;��A��.�g3ZB�ek�5W� hewئ(�T2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!D� �B���9�V��r%֌�R��������^QN�~lA�բw��Ze2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���	|e�З5�U�>�C��6�g�����t�T��?E-h��`f���sd�G}%����3fv�Cp�D�;����\���"sS<�0�zG�������&G,��G��zł)w����ۥ�Y�mK7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�;d��'�XƤ5_���H(�T�O��{Tɀ�"'��&އ�[t�Y81�d�@���G�X���.��ġ��,H�Ћ�r�H�RtV�^����ҧ|��sQ�GX�y'*��+5�4��c�L��_Yw>��������w�w:�!�`�(i3P���x�NS���U�T�C~�/b�z'hۉ)��d�7�qĉ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�@�f�smy�����B�5���U$�@p�����tA�Ɏ�A��朢֛�l����c�n�RW�A�&hH\� l���E[J��:����ڱI�̘'np>�#�=���t�T��?E-h��`f���sC>��Ӛ��S�J\7�@�f�smy╭5�k����3�]-R�\���F�`yx�>�+X�M?��y�!�`�(i3ϟ��7�4�.1p�Y,�>f5�� b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^����ҧ|��sQ�G9C�z��O�V5VM�dC��6�g��|��yp�(���z��l �>���Mb&9gUS����a$�/ϟ��7�4�4�B��Ae�,���6+�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��饭'��tA�Ɏ-՝-xC�;��|Ba���V�4|��/7*rv�n��ẹ�u`�`ÿ�����XY��\<̥�0�L�p~z�r,�)�
p�"��d���!i9�{�Jj3Ř�z��l �vPu06��K7͍���s.�֡m��z��l �M_s:Å.�g3ZB�ek�5W��x?�X�|��/7*���g�Di���0�
���b�z)�U��)���Y;e�iK!���d.���+�^n=\f�5>���ah��ol�~{�Žxjzӝ���I(͂��-��������ҧG9�:Q���ڠs^5F}���V6M��C��]��ġ��,�.���#AB��/�����>���Si��,H/��T��{B�zm&����T�3|v��Eb�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-����.�`��ai��H���9���U۸�ؽ`)[�-hn�Hlt�ٝ-@��F~*7���&�_ƃ
ᾆ�x�T�\ ���:5A��p�)��S�2�oi���:_�]4;H?�f���-A�¤�x.�Knql5R?}�b��>k�N��^��hJL��;���N�[���\��-��pQ��e��>��Օ��qvdЧ^{�j��:����
�ݚ�Н���B�1hͷ�H���9����Đ%1tSjv�!�`�(i3`)[�-hn�x�Վ��t97��EN�h�h�u+��.ᬵy���ܝi���ؼ
���$����G��s��c�!�`�(i3��jVѭ@!�`�(i3T��{B�z���b�z)le5W�F�h�j�W����Ε>�E 
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4bƗy�"c���ϰ���j�W���"�2�~�}PR�]C$�̟�1�Qטg�u2"�7 �H9-�Ԕ�k�z����\�ec[���-���d�@���G֡w�]�h��tH̾)�Z'S����7�V�Y#ѥhC�V���3������Gɟw��D��ҹnЭ:nWf���gW�6�h�g��(�K�}0Zܸ޷�d>�c�n��-��k��F*�L��!�`�(i3!�`�(i3��+�t2��������_
�u}%GP����ZLN�	���ǡ�C�a\Y����+���LQ�B����_�58���d�@���G<Ň�ć�3 �����}c��ko#�Ԯ�	\���� ���JH����8��#I�ND�s���H�V�4�(�Ҁч��ݠ�s�i�Y
�,�]�!��	Ǹ�y85���Ü�ۯm&����T��V��l/�#>6�b N>�3�eZ~��!���c�A�L'4��"�����WdM4@��hd=��&q^�`
�c��><�$��;mQ��8���/���/z*x�n;��|BE��Vˀ��e�8�ʫ��g��� |ag��6����p12���v1a{J�����X�����2�"�G�p�P�(��Iw?�d���&�Ms�����x��c�ۡ��W���\��'���Xw�j�7���4br���P[Le�/ Y�{'%s���F�p8@)y@d��4�x�Ms�����x�Y#ѥhW���\��'���Xw�j�7���4br����.J���0z�cULj� 1��Y#ѥhɠD(c!)����7���{r��'6���;8=�g��U-�e0�L���^�V��	��y ��f"䙼��"�}�k����:b����Aɺ��u`�`��c�ۡ��B�@o��[^�}� u��O���#Q�0�x3=���x�l��1:�N�*�x:��+���������i�D���K^�)��ݠ�s����M0sAo�r������-/E8�)�[���6�X;p`�g�]@n_���?3�����^�٥�@1z�+J���5���Adu�5k
��Fɴ|�O�j��O�G?X2���Y �6�ZWq�ߑ|�ҧ{�x����y���ݫ�ф���F�)k��,�:�N�*�xY��
�iCTl�������l6�Gظ0����t�%�Z?��<�ry^���"����M몴PBoTt�{#	�x�vYv�����o�|CZ�k]m��f�?ǉ�=@ E����vc]x� ��2[QvA�Xxg�H������u`�`�Y#ѥhB�@o��[^�}� u��O���#Q�0�x3=���x�l��1:�N�*�x:��+���������i�D���K^�)�y�H����M0sAo�r������-/E8�)�[���6�X;p`�g�]@n_���?3�����^�٥�@1z�+J���5���Adu�5k
��Fɴ|�O�j��O�G?X2���Y �6�ZWq�ߑ|�ҧ{�x����y���ݫ�ф���F�)k��,�:�N�*�xY��
�iCTl�������l6�Gظ0����t�%�Z?��<�ry^���"����M몴PBoTt�{#	�x�vYv����@x��r�k]m��f�?ǉ�=@ E���߹N̮�$�WdM4@�P�#��5me��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��c�.h������6���@�X6� 9��kRG���L\ ү�� �VWZ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�w܊�r%�/������0�JB�� �혅vº�w�⽒���M���o�G�m�?��˳����Z���G�dE�h�k]m��XA��v�#����G���i���ϴ�k]m���9\s�\V��	��yvѧ�_�.�����Ryr�!iD�PW����GP�d�
8�����&��`,9�H�W)�Х'���;���N���)����d���!i��nސ�ѽv1a{J��\>Pq����D�����,\��ݯbJx�nJ���yN��7��aq���N��S���nQ�rV��q�t7'�P���;^�6#9>���@]�^����C�x!�H���J��Ӊ�Z��ͺ���^E4+у��b�Bϱ����(�犽{Tɀ���S�<Ԣ��Oh��*��ġ��,���~����݁.�q�0��E|�,	㶭�
WV��	��yvѧ�_�.�a�*3���9�^>l��+t�/2����֎��ׇ��>̸*����v��6
RuB�b��~�E���W\��R�6�Z?Zaze�oY��˿^����(m�φ��<�6�@a� ��fFMqlg{y����i�q,?5qzsلx1=�I(/2]�;�6*�g�c����A(�c���_G��Hb� h�ҩ�N��	�Ȓ{A�dha#4����ʴ5��9�2�LK7͍��|��W&":��=����t/�����sc�̆�!Y�X��9K`lk��`dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩΗ�nސ�ѽv1a{J��;�6*`lk��`�������iA'R�	�$(�G�����Q����$�!b���9�}4Ŀ�ЈH�����b�'Beͧ��&�~LI���p��9�2�L�Ɔ �����O�����O�ALQ�'�i�*�쳝]Ņ�*"���"fĉ>99��A0ok�����F��O�\E�W��4b��os�鮊��~TX��MUǪ�^ZE�S�8w�b��Shw��k]m���I����~u�Ɔ �����O�����;���=L�וc��f���u*Z�������5ʦ�i;��#��F�r�f�tm�;����Ɔ ���.�&�?���DKY���k]m��F���d H@48բ�z�וc��f���u*Z����9mh��n,2$����;^�6#9>���@]�l�uV�2j��=��
��d���m��+�Z����y�=��X�t�iZ]XF�hx��G��N����p$��<
DN͗&8�,�nU�gF�r�f�t���MK�L��.��֞�������i�4��%�;��g��cH�wA�?�D�g��ۤ���ֻ���~��a[/������N�� �ȳT�_�O�0Pa!�����V�`�4G&��z�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cUL#������b�'BeWh4:z�]MD�wP�/�wK��=�C�b�'BeXxg�H���M? D����j��=��
�lo3��$����'HY-��
�C�+6�1����K9
��ЅT�,\ަ�It'N�����N����p$��<
DN͗&8�,�nU�gF�r�f�ts4��u�($Q
ˋ!E\1�1�ҕ-����s�;�9�����:�.�9���T�I����1�kCW�O a�Ɔ ����û�/����q�����@�yc
׬sQ�9�&��*���j�ׇӭ��ss2����
)\Y�����'u���ɿJ�ׇӭ���W�"�Ů7��B����3�=������Fz��2*Q=F���q/���<��"F��j�u(k�ɩ4@Q�/����Fz�k/�z�xEQ���*[UxG���Fz����ꀍ�˺�Q���8X�˞�DG��9��稕�a�/!O�8X�˞�DG �@��&}��s�H��rs�i��='̹Z�;�C�x!�H��dm��u�ׇӭ��p�n��.!ū�ez��k]m��)�P�ap�>f��+�42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN%ڤ L���V��m[=��slc�����T!�P�謃@9$7��T�9=3�gK��@g2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�&�؛�$dkǔ�ˌ�1��\��L�FZ�1����ǲ]��=�w������K���'�Y�Y`$�E�.1p�Y,�-��h����F����Fu^��0�M�&�^������t�T��?E-h��`f���sd�G}%����3fv�Cp�D�;����\���"sS<�0�zG�������&G,��G��z�T�B�X
���*(H=�ƍ2���l�����g�Z��3��a���!@�f")u��r��܌;���'����u��r�妷��ҧ|���|��vz �δ��NEP�B�����n�(��&������ҧ|���|��pr�<:\��
�
��(am�b3�D�4���܂W�/�#+*f|���|��pr�<:\��
�
��(8�Z5	Aݨg��U-�e2�B���7.�`��ai��NEP�B+�,�=[�le5W�F�h��
�
��(���>05H~fĉ>99��A0ok�����F��O�\E�W��4bƗy�"c���ϰ��턭
�
��(�o��!���=b��uǓk`���)9`���M#��y>'MM귈nIg�R�5��/dV�ļަ��P���]6����(����c�n�R�HM���#g�8����f���-A�¤�x.�Knq���;W��ZLN�	���M�X�FG�p�P�➁q��H�g 6ͥk�0�=<MW�-}�	mp,��_А#�<om���ug�RM�;��|Bq�D�7�j����tL�M����
���R8�+��@-�-'͏�������x{�~�WR�7h�,b0V�u�Q�ݚ�Н��
�I�>y!�`�(i3��i�\�{q����W�Ty��5!�`�(i3�gCu(o?C!�`�(i3LZR���[������2������}F�G���d2������}��s�5e��g��cH�wA�?�ۖ0����[� �GR��shbvk~�#x ��M��.ᬵy��ݼ?����DY~�y����o)�T*�c��n�da�ۣ���(�犽{Tɀ�$����nQ�rV,?����)�{6�U��ΡKCh��(	�G��^����K�7����&Y��V�ǣ©��$��:�e�hfH'��!�i����VZDf�?ǉ�=�O�G?X2�K��2WI'�=��yp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���m�
��,!q�\E��0D������'���Xw�j�7���Ɔ ���9/�^Â�wӨj]h����dЕi�����,��%�N�dТ���S֜���,�ǰ�98#.�Ƌ�Z{oBQ��;��O�"�Yi���t�E��j�AkUx���6�|����CԀ"<�h^�hvl��9�h �=������-�S�h �=�*�a"4̥�0�L�p~z�r,��:fۇ�0�=<MW�-}�	mp,��_А#�<om���Ϻ� ��H����8�(����������cɧ �GR��shbvk~�#x ��M��.ᬵy�����	��u a⣃_B�h���Q�kUx���6hnp7�=Z鎬�������(���'�jh�,o�"ɑ�聾.�g3Z�Ǵݵ�������� �a���GE�A�'G���f݄pB��j��=b��u�_3GH�F���E���b��y>'MM귈nIg�R�5��/dV�ļަ��P���]6����(����c�n�R�HM���#g�`Bu�������}>p~z�r,�+�/��f���-A�¤�x.�Knq���;W��ZLN�	���M�X�FG�p�P�➁q��H�g 6ͥk�0�=<MW�-}�	mp,��_А#�<om���ug�RM�;��|Bq�D�7�j����tL�M������>r���+��@-�-'͏�������x{�~�WR�7h�,b0V�u�Q�ݚ�Н��
�I�>y!�`�(i3��i�\�{q����W�Ty��5!�`�(i3�gCu(o?C!�`�(i3LZR���[������2������}F�G���d2������}��s�5e��g��cH�wA�?�p�p�{V'��kd.Cf����+9��lE딧 �GR��shbvk~�#x ��M��.ᬵy��ݼ?����DY~�y����o)�T*�c��n�da�ۣ���(�犽{Tɀ�$����nQ�rV,?�����k��M���'abW�5�}�]��ϵ��t�pu:�]f�?ǉ�=�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��W�"�Ů7�6��,�ݜt���,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ:��IK��<[�л���7M+э4��Y�{'%s��jb�ܳ�/�����b>I�Wkxf�?ǉ�=D�wP�/�w���bc��U�d�#�by��W��;_��8W�w��fD)IA����Cj����tLB�'�4V�������� �a���GE���T��>f�l0 ��J��9j.�l>'�o��&L�/<�t��Cn��P)��	�+�`g�]@n_���?3+��y(��'{}yw~�귈nIg�R�5��/dV�L�溥����v�8:ۛ@W:���#���F��*{�욋�Օ��qvdЧ^{�j)�]�T��z�**ߜ�*�l8�b(������l__��E� )�&,�W�8"M�5�O�%E#Pڗ����7���T��>̷_��yC��S8�vV�y��F�k]m�������%�w�R���y �+�5�?+�T��ˬ8��� �r-��M�s�����%8&�d�I�_#�	�Zz/3>��-��k�5��05N)hiW�U����҉�p��P���x�a[M��1�:�Ω�����|"����T�N�R�7h�,b0V�u�Q��M�=�@���k��!�`�(i3��4��#o�;-;*�7����E�����-/E8�)�[���6�X;p`��ļަ��P�5��/dV~����G귈nIg�R�5��/dV��H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	�螎X�zgz�'�̗���������D�ڐD�f�.���ژ��V
�E.Q�,��SOV��̺g�z�)%/������Ó�U kuB�b�E8�9������ցe���ɯ;�{d��L������
��3x�,� ΡKCh��(	�G��^����K�7����&Y��V�ǣ©���W�"�Ů7��B����3�=���jo�����<o���D�噸��\i�s�h?��dv��oTN֢&@��&�M�g����H��bf�?ǉ�=���ꀍ�˺�Q���f�?ǉ�=&��s���qz�Gb��P��2��}��CϾH�)�]�!��	Ǹ�y85��J��ꅙ��uF��t�{#	�x����dЕi�����,�S=���L�X�{Yr�<�؝�Z�^lj��b>|�~n�~/�k��?΀�(4��AYp<#��v�5M/~֔��p�;v�[�I�?g�f&:��r-,ب���H��ϸ��#|S������3[�u8�U��֜��3!�`�(i3�kޮ��n���㬺j;��q,$Q
ˋ!E\1�1�ҕ-��'{}yw~�귈nIg�R!�ZV)}f�~����G귈nIg�R�5��/dV��� �"�W�A�&hH\r��ي�2f���-A�¤�x.�Knq	6�q�i�d�<om���!$��x5H����8�裖M���"�c���ژ��V
�E.Q�,��SOV��̺g�z�)%/������Ó�U kuB�b�E8�9������ցe���ɯ;�{d��L������
��3x�,� ΡKCh��(	�G��^����K�7����&Y��V�ǣ©���W�"�Ů7��B����3�=���jo�����<o���D�噸��\i�s�h?��dv��oTN֢&@��&�M�g����H��bf�?ǉ�=���ꀍ�˺�Q���f�?ǉ�=&��s���qz�Gb��P��2��}��CϾH�)�]�!��	Ǹ�y85��J���K�+���w��@IAE�{k�h�+�>��y��j����tL'�xx0{�|ag��6���6*E�}���2$e�i7N�_�z*K��I4��欱���j����Eo(d�J��:����/�M�í��{_xGSnǀ��+Z}�E+8�D�}����Tf���-A�¤�x.�Knq	6�q�i�d�<om��إ�E��c���$1&O�#�-�p�~�Y����.����j��k��?��,\���yr�/ӶWȶ���/�Z�k�ʆ-�(i�pY%���m��3��p���H����HRCJ��<om���o�p��F��0,5 .�U%{.�V#?p�&���A��id I����*y}e��=2�������4}�5:����97��ENҨ�ᙨ�vuƇgv)���N�N�q*�CO��0�=<MW�-}�	mp����"���;���N���q���4!����~JC�[��~f�� l����jA��L�L�溥����v�8:hJ�tV�nQ�rV~��s�N�$²�ؗ$_\���.7
��l^U�L�E��w*�8.����6��}Dq�f�˥�'ܤ",����=�˨6�o8:4�I���c�90B3v�A��d=��¾ȼ!�`�(i3�'ž1�|�'����u��r��L��@�a��Hb�2�Ǐ�iA'R�	��)���Ҟ������'���Xw�j�7�����P�|T��D�?��/��j����?zk�8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt> #6��r��������]�YW�Z\PН�l�����=̞��>�h�5,Wlr�r%)cA�1#V���<e��ȅ*Ghy�`�w��v1a{J��]V9��WҞ������'���Xw�j�7�����P�|T��D�?��/��j����?zk�8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt�j��F=W���}���i���>8I�p_�Gt�7A�;�֋`NY~�y����u{ᵿ����ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��=�O�-v�*�Va�irv�A�
^^3�V�C��k���a�K�v�A�
^^3�V�C��k���T�7:-�w���+_�mS8<�n�ݚ�Н�F<�����R��1tSjv�!�`�(i3���$Q�@=��X��/�-oRCGtKż���b�氦�=��X��/�-oRCGtKż��9*�����!�`�(i3m�ľZ��*!�`�(i3m�����Gd��}U؄�k]m�����m;
h�����B]�PZ鎬�������(����,F(dA�F�u�����j W'G�ݚ�Н��������;�P�t�5!�`�(i3��p`-�F/͘6��q��kUx���6��~�^AԢ�a\蟹D��wX��n���㬺Q̹Z��u��r��!�`�(i3�S�y"�J���.!G@��Hb�2�Ǐ�iA'R�	��)��޾���gf�� l��}I�?d�G5V������yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a�*&\�{I�ٝ�z*���q3+Ԣ�0�=<MW�-}�	mp����"���;���N���q���4!����~4�����ݚ�Н�!�`�(i3v���,Ͽ�2[QvA�ͧ��&�~L~l�d����!���c�A�L'�ɻ������+��<�ao����O����8Q����ze�x�T�ݚ�Н�
�:qEp'{w#/ B!�`�(i3��k�C�-�<�ao����O����8Q������51�X�c�rs�i�}�O��L��_
�uk*����S�~���e�)qP@L0��U���(�犽{Tɀ�$����J�	�LÆ��S1�c������b5?H" 1����>E�%��*d��:=�;�մN���_�Gt�7A�;�֋`NY~�y����u{ᵿ����ݚ�Н�
�:qEp�;�P�t�5!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��W?�;��5��S*#���{�6�EZi˒ow�R���y>��yС��#x���.1�	;�IV��o5]�$˹�+�P�ф�?�s�5@䯁j]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M��b�p����ī�����vM�)���\���F�`yx�>�+X�M?��y�!�`�(i3v�A�
^^3�V�C��k�&�c���R�NTgccv%��v��!�`�(i3v�A�
^^3�V�C��k�&�c��������	p'��$�\%e��}Dq�f���9��稕/Tu���Ŝ��%ٿ���H�w�l�ß�
s��ƍ2���l�N
����\� C&����q��Z��V�X8�9a �<�5Ɂ7)P<�ܓ�Y��+�t2�����dz����NR�p��@���|2~�|��� �ҋ�;��}Dq�f�dl��[�����{�6�*F=ॵ��@x��e�d�$7 �ҋ�;��}Dq�f�dl��[�����{�6��q��Z��l:qvB�%��v��՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r�剅�%>�rGWfי�b����{�6�9\�B^6�/.�<�����&aD�4�X�X�>c�.A�(��cS�c�X�X�>c�.A���BO�#��}Dq�f��6[��u����@~H�k����`T�]b ����ji���&aD�4�X�X�>c�.A���d���T���@~H��k]m��/r����1�ߤ�:C
#!�`�(i3v�A�
^^3�V�C��k�&�c���f�s栿o�x�`�8�Gl�x����b�'Be��/=��v�A�
^^3�V�C��k�HvL)��x�l�����}Dq�f�N
����\� C&����q��Z��V�X8�9a �<�5Ɂ7��C�=�g4�B��2�k1�h�H��*�*���\� C&����q��Z����/ǭ�� ��j���ݚ�Н��f���My���O��H�ߝ�;�K��CL�УΛ
V��q������5*g]�H�X��%�CV߯_-��+�t2�����dz����NR�p��@���|2~�|�����:l��0�5G,��Gc#�ѿKM'4˒���dz����NR�p�+yG_��\�����a�)�1�׀�<�6�Q==z!
���-�F�i��|�Uk�rDp!!v*!���K�5OoL!���}/
;$�Z��"�Y�<�SЮ!�`�(i3dl��[�����{�6�*F=ॵ��@x��e�d�$7/̉�#��_�X�X�>M�a���;}`O�kХf�Q���V�C��k����?dq���z����7ir	� EG���͵u����p�����+X��FJ���-�����ND��_�W�.��;�#5�UWF�g���On�T.M!�`�(i3R��ak����`T1�h�H��*������AZ�,��#�2
��e���.��;�#;Y���@+���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�~(����W������Ȃ�`u�'���Y^y�*ܦ��&Y��V�����^������=�˨6�o8:4�I���c�90B3v�A��{y����i�q,?5qzsلx1=t�0��@�E$�I�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�u����p��8��V\�J#�	g���=<�6>e��0�U+�qbp@�!�`�(i3zk����G7```+��BM"�n��>�my$�N��o�/���;��+�t2�����V���V�%�1⢄1@aw5b_X�XV�b�z'hۉ)��d�7�qĘV�52SG�U��@at3Y��P4v��*����E�g�������(ӈ���m�r���������y+��
 A�O֦�w�#d�R�NTgccv��nF���<�W�.�P�	��
�Q�}uD�*';;���41IL����֟D��m#?dN�<@Iv��nt=:��:5A��pG� �l
s����9�~��� �������Z;P��b+}y[�V�52SG�U��@atA�ᴽ�����_�q9+t�}�ݚ�Н�v���,Ͽ�2[QvA�%ρ��r�/ ���we��0�U+�qbp@�!�`�(i3�@��A���k]m��>�,��,� n��>�my$�N��o�/���;�q�9�ͭhy�`�w��v1a{J���A�qx����E2b�z'hۉ)��d�7�q�L��@�a��FD>�v��Pn<���*:k(v�E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*�Va�irv�A�
^^3�V�C��k�&�c��������	p'G��Hb� h�ҩ�7�wtMM���j�=Nb����d�3��[(��}�%Dܭ5�4-+EsҤyM�d�X'�i�*ڶ�UKs,��l�?�C�g�k`���)م�_ҩn!�`�(i3zk����G7```+��BM"�'�Z��ƾU��@at�f�6l�}sf�e�}s�dKa���^�uPϿ.U�d�#�b��97y��!�`�(i3�?�:>ɡ?�s^�PD�9������MV�,o�����&G!�`�(i3/w1z��ӊx�D�Re|����x����,����_
�u�2��Y�f��y	����F��،!|�α+
�:qEp'{w#/ B!�`�(i3o� c �R�%1���%��K��>P��}�%Dܭ�ߦ?�~F��C~/*�xK���&T!�`�(i3���F��O��ݚ�Н�G� �l
s����9�~��� ������ESҩzk�����>�P,љIX�o%. *.�ݚ�Н��e�<Q���c�ۡ��ZiC����I����~uAԢ�a\�ۯ���@Z�2[QvA�&u�)m��J�e��RWL��@�a��Hb�2�Ǐ��Pn<���*:k(v�/g��6��c�ۡ��ZiC�����}Dq�f���Ě�����}Dq�f�܌;���d��-��!i��$>�cQ׆��p0~�5�HRoP��e��I�߷�c/��-����!�`�(i3����6`X�/m>8Φ�ck��x��ɪ�����:~�Y����.��������h�4��=y����͘6��q��kUx���6{��.���ݚ�Н�G� �l
s�M��K��'�,LF���ji����V��G �pȌ���]���E:�qL��n��p��b�Bϱ�fePh��������9��}Dq�f�L��/\��=2���H��̣��R�)�	8k��.ͥ�H�RtV�^��.J7h����ly�P�r��n�Ŀht�2�q㬑�,\��ݝۺ���r��������]�Y�_�H��!�`�(i3�����!�`�(i3/w1z��ӊx�D�Re���x��O ������:~�Y���Wql���8z8�t�RL��}Dq�f�HN��R��bP�63Z�t�V�52SG�U��@atA�ᴽ�����_�
w�	������9�~�nI��Y��!�@�VҒm�L��@�a��FD>�v��Pn<���@���(9[���G�������+��+�g�>U�#!��&vY��;��q�9�ͭ�n�Jt�g�v1a{J���A�q�3�4�f��+�g�>U6���z�S�:5A��p$f��_Ub����B�)�{6�U�����F��O�}�	76�&�φ��<�6��o�u�/��Rlj���H����t~�vE�s?�s^�PD�9����%�줝v)ڥ����Ⱦzk����G7```+��BM"��O�&��̏�c�ۡ��ZiC����~eWSQl�\� C&����q��Z��V�X8�9aO�˰�]q���X��O�m�4VGG� �l
s����9�~�nI��Y��!��N��rJ��Ű#����=2��b����d��i�8�����W�W[��m�U��k/�ț��OP�˟D��_�W�.��;�#��f��w�f� .):ާ���虾�b+}y[dl��[�����{�6��q��Z������5�r�M�{�|L��!ߩ��`4%�fZF�Gck��x����,��
e����j�=Nb����d��i�8�%m�Y$� 1<F� �����C�D��K�֢��s�Kȓ�FG����3�4�f��<�ao���CC���ˊ�ki�3zk�����>�P,љI�D��|�|-��4��C�;_�b�z'hۉ)��d�7�q���}F�*B��F�f�J���1��]/g��6�Y#ѥhUM�;Se<���j�R��=2���H��̣��h��b����wl53�e�'{w#/ B!�`�(i3!�`�(i3!�`�(i3�,\����Z:@��@W���}���i���R��|}&���Tum��T˥�'ܤ",����^�� �YW;C����bi3�I�߷�c/횆����X�X�񳱅���^����zlv�]w4W�'{w#/ B!�`�(i3!�`�(i3!�`�(i3�{_8�Y��=�}�Vݨ-n���n�v�ĺ�֦�w�#d�m��u/�Οt�,�NL}�="��x8I��Ig"�R�o� c �R�%1���%HIm�T���x�bG�Uew���m����x��O ��f�����&Sq�aL����֟D�ʥҔFܽ���ly�P�r��n�Ŀh9�-�wQ�ؾ#(�[�(D��_�W���$� 8C��D9�C3x�В&=�y�q}��5,�����t�iZ]XF�hx��G��!�`�(i3U��֜��3!�`�(i3X�PC!v�@[�JJ1��P�M��,���9^-���.��֞�������i�_o�dZ � �GR��shbvk~�#xǩ"�4s2nQ�rVA�H��%��SFU� �hΡKCh��(	�G��^����K�7����&Y��V�ǣ©��$��:�e�hfH'��!�i����VZDf�?ǉ�=�O�G?X2�K��2WI'�=��yp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���m�
��,!q�\E��0D������'���Xw�j�7���ڹ�)�u="��x8I���A�-!�`�(i3@ E���߲	[F42��c�ۡ�����Ƭ��,@�n���r�XB�a���?7��au��at�kZ+��T�����D3��־���1PM�^-q�x�l��1:�N�*�x¥������]n��-��%{.�V#?p�&���A	{K�tU�P!�`�(i3�gCu(o?C!�`�(i3zR��_��m��3��p���H����Q#�?���;���Nxk�~̔=Z!�`�(i3^P��:w0I� X�1�;LV^Š�r��Lo�_!�`�(i3�2*Q=F�k�mD#V��A��`-2Y��kک�x����y���ݫ�ф���F�)�_�������� "5�]�B�'��a�F�,�U6�Q�L���/��@��:$����z�����	�;�ݚ�Н���"����M몴PBoT�ݚ�Н���_(x��`g�%Y��̗0z�cUL��s@OĪkew���m����x��O hH�
$;�?V��j�c�;J�*%n��@��A���k]m�����2�¤Ƕ�W�I&!y'}�}c��ko#�W��xS�v���,Ͽ�2[QvA�ͧ��&�~L]���E:�qL��n��p��b�Bϱ�fePh������w9���e�<Q��Y#ѥh��Ů@�	����W�W}c��ko#��J��Ӊ��@�#��ErS�b�8Z�AԢ�a\��!��a�'�A�Y��|s����"h�ؾ#(�[�(��Cn��%�<'L�+��T�����D3��־���1PM�^-q�x�l��1:�N�*�x¥������]n��-��%{.�V#?p�&���A	{K�tU�P!�`�(i3�gCu(o?C!�`�(i3y�Z�;���>0�1ۍ�h �=�f�?ǉ�=��'abW�5�}�]��ϵ��t�pu:�]f�?ǉ�=�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��W�"�Ů7�6��,�ݜt���,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ:��IK��<[�л���7�~@M��@�Hb�2�Ǐ�t*����B7Ԅ��{k�h�+�0��NZ�Hb�2�Ǐ��t���	�%�% ��5���"�@��A�ی:�Gɩ��I�?g�f&:��r-,ب���H������%kR��������֢&@��&��x��&^�B�wj$g�X;p`�r��������]�YY'K�"M�,�zg��p�r�X�<\�!�`�(i3�����
L�c�n�R�V�E�-�9�ݚ�Н�ss2����
)\Y�����'u���ɿJ��ݚ�Н��W�"�Ů7��B����3�=���!�`�(i3�2*Q=F���q/���<�����7
�e����kn4@Q�/�!�`�(i3k/�z�xEQ���*[UxG!�`�(i3���ꀍ�˺�Q���f�?ǉ�=��9��稕�a�/!O�f�?ǉ�= �@��&}��{� �Q ���3���Ι��Ȣy�!f�?ǉ�=D�wP�/�w�!�v���3���΂�l/�Q�e����M<��}�u�?�d���&�/�M�í��'���H��1%��D,6j�"Hsη�m\
�NK��v�nJZ#Je޶^2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�![�,�ᖠ��I�v�o2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�|�)՜�4����;qX�qp�c� xG.�w��G�}CL+�J���,�)HVi�pz��AY���Z�@���v��d�-td'�I1L�S�Xr&ߜ����nPB���׭'wH^��Ƨ�0͜��!?@K���୩���&�K�VF�T֣[\5Cw�Hm�̶^�+3��F-|S5�g��L�*� )�\�~xy���T�}ɻY~�y�����[�T���Ӫ!�J��:����Qw�$��Z��/�dW�<龈��ơlП���V03Y��9�`�I��W����Ľ��M�ȅõ����(�x�HM���#g�s�
�`�I��W�^��D����jVѭ@!�`�(i3!�`�(i3!�`�(i3S`�@���;_��8W�w��fD���4s1�L9�_�mEn��8�g�^[�q�eʣ͜��.�4�Bg �A�o�Ղ�f��T0	�]T��Fn{�^l�tċ^9t���G���U��C!]cq���<�&i)$|�&��YTi�#�~�H:$�Qo�4L�⨴��[0V4�*��:&���#��)�824F���ZٱNNu�A���r!B�8��`ɂw���:.�\����@�����`�#}�{�u`nWM����l�Oc�d���]�c�$ͯ��L9�_�mE3��<t���r�Ŏ�]ΟQ��ǺΕR��ӟ-�ЕS�#m,�t��gJB��#U#��F�	�l�V帐:ŧq�J��:����Qw�$��Z��/�dW�<龈��ơlП���V03Y��9�`�I��W����Ľ��M�ȅõ����(�x�HM���#gO"J#]"+G��~�I��T+Ĺ����ġ��,
�����F��]#��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3پ[���-��Z?�6j�"Hs!�pL_�g��L�*� )�\�~xy�������4�-���G$��S��n��¤�x%��u%�RA�8�>r&�G�p�P�CX�p1����6cox�%�/��Z>L�0������H!�z�l��d���!i���jSA n2ϒ���=��pȠ��ղ]��G��-y�� ����i9vo��ob$fAԢ�a\�\���V#��p~z�r,�ܯ�kC�4��]#��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3پ[���-��Z?�6j�"Hs!�pL_�g��L�*� )�\�~xy:jT��J���9��稕/Tu�����_&�����d���V�M�{�|L����5m��Y�j�`M4��c�����:/��N��׮	��48ܼ�P���6�5>EZU2��53��O��h$)��� �GR��shbvk~�#x ��M��.ᬵy��b��k�|��n쯎+�ܼ�P����JhF�Ԯї9gP�U,�2������}��6�L�-).^QQ#j�o�������԰����H-�-�o%�_�*�@W!�`�(i3!�`�(i3!�`�(i3!�`�(i3��b+}y[v�A�
^^3�V�C��k�HvL)��&d��]�^���H> �V03Y��9�`�I��WF�\F�l9Z��b�Bϱ����(��g.Cf���Ϲ��,䮰�_�B&��p�+9��lE딧 �GR��shbvk~�#x ��M��.ᬵy��ݼ?����DY~�y����o)�T*�c����g\�,T:5�����2������}Ov�xIBB[|��;�ċ�lʥԊϭ�Ī��$b4i� ����i9v��խd}���![<b/�>Ac�'{}yw~�귈nIg�R�5��/dV��s�;�9�����:�.�B7�-�6!�`�(i3!�`�(i3!�`�(i3!�`�(i3��b+}y[v�A�
^^3�V�C��k�HvL)���g��L*^���H> �V03Y��9�`�I��WF�\F�l9Z��b�Bϱ����(��g.Cf���Ϲ��,䮰�_�B&��p��ey��qE0�n쯎+�ܼ�P���(�K�g���yN��7��aq��G�n���t�;���NI	��y7DT?�R��n}�����H�i
�J���̥�0�L�p~z�r,n}_��嗍d&�.�_�L[� �h�����T)#�y�ö�7�-).^QQ#j�o�������԰�W����V'��kd.Cf����)Y����2�g�]@n_���?3B��A���!�`�(i3!�`�(i3!�`�(i3!�`�(i3`/v�!!]�L�����B��2�k1�h�H��*��iI������x������p'7T\� C&����q��Z���2%�ɛ'���$� ���u�,4	M����ge��L�����B��2�k1�h�H��*����p���x������p'7T\� C&����q��Z���2%�ɛ'�F7�Gh��r��C�M����ge�=���r�%G�Y#ѥh�g8V#��4֡\�`!|��{�7{�2z����!Cu�>(���] 9�X� U�X����d���!iZ�,��#�2
��e�������m[�LEE�S��-��h��ڥ����Ⱦq���3��`��R�`�mQ�x�z�oi���:�&2u/H���(�犽{Tɀ�$����nQ�rV���#����}�YЦJ%I!Cu�>(���] 9��/��ʲ��n2^���;_��8W�w��fD�@��A��2��� �ЁV��vD�����m[�EBS<u����3���΢#�7�
�k
��d��6�����m[�~m���Z���n����o/i�\	t��H��[k��q��־pT��sP�/Tu����W`GU�!i&G�\��u��6��+(c�q9+t�}�t����M~V��	��y'��j���+�g�>U�� t��{��X��"��ҩ�	rGf��x��9	4��t�f!�`�(i3J�a$�Y ^���H> �?N\z��И���|�bo��ob$fAԢ�a\�Zx�.����#�喵K��zd���|�b��խd�g��;�!�`�(i3!�`�(i3�>d�g�K�9;��ˉC�G����]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7��k���;\�Dj#.�\���F�`yx�>�+X�M?��yЛ���a���2�6�d�f%��v�ڕd�tuѭE��ȷ��%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3+���G���9�+��N�=	�N��!�`�(i3#� �,W�j�o�u����-Q�OPHN��R��bP�63Z�t�5ߧE4��Fr��j��k���;V�
pFV��ۄI��K��I��gs7ߐ)�~ң>0�1ۍ�h �=��Y��"��5�O�%E#P�Ͱ�Ǭ�j��e���W������)<��U��)���Y;e�iK!���d.O.C�U��B��-����A�;�����\��]8��	�����;c�~�r$ɓǃl[�Ƶ�1tSjv�.��J���nz�����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv��/��@��t��ܜ�[�E��y���'%������e.��>�g��U-�er�.�j {:fh�3�:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��o�.�u:u����<�x���ަЅ.�g3Zꢯ�wv���`	HX'�NxPr[-]�e���?ͧg.~�-%H��s�;�9�����:�.U��~��� a⣃_B����ѥ�)t��ܜ�[�dN�<@Iv��;z�����{:fh�3�'�֝�p6j�"Hs�c)�W]��P�),�w���� y���t�T��?E-h��`f���sd�G}%����3fX�?���'��>��ԑ�%xjzӝ���I(͂��-����N
����e���b�!�`�(i3!�`�(i3J�a$�Y )P<�ܓ�Y��ɕ�eYl�x����b�'Be�s�r��<�!�`�(i3��nF���<�W�.�P�	��
�Q�}��9��稕/Tu�����_&�����-陹��J�a$�Y dN�<@Iv��nt=:��:5A��p&aD�4�X�X�>c�.A��I�JZ����;q�{_8�Y��=�}�Vݨ��}Dq�f�q���3��`��R�`�mQ�x�z�oi���:�AS#��]�,\�����O��x§0�=<MW�-}�	mp,��_А#�<om��L�'Ҩ肋@�Af8�ٕ��(�W�!Ċ&���X�G[�x���01�m+�D8t�R!ME�D��_�W�.��;�#��&�qҸ�2Mz`���^E4+у��b�Bϱ��L�溥����v�8:ۛ@W:���#���F�Q+o�>u����p�����+X��FJ���-],��%s��(_w�i�<�<j��.#�#�-�p�@�Af8�ٕ��(�Wl N��~�!�`�(i3/ ���we��0�U+�qbp@��#�-�p�@�Af8�ٕ��(�W.�pڃY!�`�(i3/ ���we��0�U+�qbp@�</Sn��/Tu����W`GU�!i&G�\��uG$�ء�/ ���we��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3V@���gx2!�`�(i3!�`�(i3�	��*��)-�8�ήu��}Dq�f���9��稕/Tu�����_&���L��)%�4Wfי�b��}!D̅��}���wWfי�b��}!D̅����A���r�>p�{C��Nq~o@&aD�4�X�X�>c�.A�����WՉ��%>�rGWfי�b��}!D̅����<!GO#B�t�x���@~H��k]m��E7�y�PjNh���W<˥�'ܤ",��E� ���_w�?��g��U-�e�����1l�x����b�'Be��
�����V+���]��ɕ�eYl�x����b�'Be
��e,�U�s
ƺQ׆��p0�Ĝ(�IyIR�%r?�	rWfי�b��}!D̅��t/)����ݵ�Q�n��T�\ �͉ק��l����@~H��k]m���V'��KchL<D��`0`���*17�wtMM�0�5G,��Gc#�T�Ed�	��*��\� C&����q��Z��NH��\-{@�Af8�ٕ��(�W�W���+@ܑ��y���8���/�>�h��fLD��_�W�.��;�#$@�s>�
՜�}Dq�f��L�����B��2�k1�h�H��*���ެ��u����p�����+X��FJ���-�����ND��_�W�.��;�#5�UWF�g�9gUS����a$�/q���3��`��R�`�mQ�x�z��1�K�!�/��@��A���3A�n�+�sQ}b`������	�%1AZ�,��#�2
��e�������m[�P�j�OD;�R��ak����`T�ҩ�	r^A�Y���b�������Cҷ��eHy�\D������{�6�*F=ॵ��@x����W�HN��R��bP�63Z�t܌;���d��-��!i��$>�cQ׆��p0�Ĝ(�IyI�I�CPWfי�b��}!D̅����<!GO#՝�]�k����geE�vx���ƚPyeP��m��'����C;����Hu�S��%� <9[�Z�Wm���Xb�z�Ou��y�:n�%\��Gݫ,��G�.Y@NJׯF��G?Ґ80�)�n8q����JA����2����:&�)m���l��֘�^��A�l��><�e�BH1iV�x��8<�@�Af8�ٕ��(�W�!Ċ&���X�G[�*����21tSjv���+�t2�����dz����NR�p�'q�-��nEg�N>Z�s���Wwq���3��`��R�`�mQ�x�z�oi���:4#��^x���ݚ�Н����F��O��;b�-�2��;�P�t�5�H�����Yu���*Y��b"Wfי�b��}!D̅��t/)����(��cS�c�X�X�>c�.A�L]�f��e��������Oݥ��{)�h �=�$��bY\���ZAL�:y�g��K��7�I�$Q�ϐ �S���pj; �B�o�+�m
Og:Ba=�u��Y'G�vw�B��qbb��fddf�ݲ�UC֬g'�J|���������k{s�^,ysA�U�y��6��3fU����O���X#��cA;�jmT�#u����p�����+X��FJ���-],��%s���fcŘ��v��ONH!�`�(i3�L�����B��2�k1�h�H��*F7	G�<�*��s��ꮂ��}�%DܭD��_�W�.��;�#��&�qҸ�2Mz`����G�x )HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�2oY��.��x�13�K��oNYzZF����9��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7���z�G�	S�uimK������t�r$ɓǃl[�Ƶ�1tSjv� �#0xg�`�I��Wn��>�my$�N��o�/���;����������zՠ�����˦G�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�>��:J�E�<����i"����*ȑs��,:&�^��,Q����-����!�`�(i3R�c4!`��Bf���Q١Ӿ�$���l�K�F���m¡HN��R��bP�63Z�ta�F�������Y���D��3��bt�u�&��F�ߏ��D厺��+�̟�1��$!��8�ZLN�	��l��Z�C�H�RtV�^>�Q�c6�����-ќv�Y_�R��D厺��+���l�K�>��������w�w:�!�`�(i3gJy��8���O?����'DV���b�z'hۉ)��d�7�qĉ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j���z�G�	S�uimK�(�ޞ��]i�ţ��t,�� .6�o8:4�I���c�90��G��6�iI9�o«IX0F�M��ŊPTWo9�����j���A(�c���_G��Hb� h�ҩ�ʬw�S���q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�ʬw�S��ht��p���j��8�u��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���]i�ţ���Al+�H�R�7ʌ�J����φ��<�6�@a� ��fFMqlg{y����i�q,?5q�+�#4��F��8M���"sS<�0�zG�������&G?V��j�c��׽��dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ��)��S�2�oi���:_�]4;H?�f���-A�¤�x.�Knql5R?}�b��>k�N��^��hJL��;���N���l_�c�u��r���2��}�����3R�� ,��rQ͒������ݚ�Н���jVѭ@!�`�(i3�4�	��3|v��Eb�z'hۉ)��d�7�qĉ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�@�f�smyP�@Ե5����EO��]C�1�kU�i������ ���JH����8��#I�ND�s���H�V�n8�A�A���p��b��!���?t��my$�N��o�/���;w�R���y����<�..�4���R@�6���*��ˌ�t3�{E��'Z*)�?�R��nj��P_Q����t�h��W+��W�v,���cL�Ec'�\Y-φ��<�6�@a� ��fFMqlg�2N��n��W�Q��a�U��@�fћ7��'�b���b�Bϱ���w�K���1`��vߜ�*�l8�b(������#oMZ�n��[��{_8�Y��=�}�Vݨ��}Dq�f� ��b�FP&�YN
��)ej{�y���q��T�ٮ|�,
���A�;�֋`NY~�y����u{ᵿ�����"X��[�������q(����b�z'hۉ)��d�7�qħ2N��n��E��������Z��o���i�#Ѻ'���Xw�j�7���kv޶Gla��Mp�g��U-�ei�X'H�;C@�����{_8�Y��=�}�Vݨݾ�9J�ciI9�o«IX0F�M��ŊPTWo9����'��Q��r$ɓǃl[�Ƶ�1tSjv�џ�3~�l"U��@�fћ������K7͍��|��W&":�ݚ�Н��YN
��)ej{�y���l|�*"k���(ӈ���m�r����(1l�jG���Z��oYTZ�@�K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv��B�'��a���p��b��x��f���!���c�A�L'��B9[���a����}Dq�f�hs�����n��0�5	x�qr�~����p��b���1�ͺ'�!�`�(i3�%�r���°��Yzw�x��w�����&����!�$�Rľ%�� �GR��shbvk~�#x��	���1tSjv�!�`�(i3͝�����|VO�⅘����-a������aGl�6 y2��R�՝� s�#t��ۻz���Yu��^��.�mZ����������yN��7��aq��zW�&��F�u��r��!�`�(i3���e�T�%�td7���{_8�Y��=�}�Vݨ��}Dq�f�;�jmT�#�YN
��)e
Q��fh�5,Wlr�r%)cA/�r�]/2�ݚ�Н��B�'��a�S���%���aH(���{S���%��jYȺ8�8�!�`�(i3�	��x��ݚ�Н��B�'��a�S���%��V�O��%��e��0�U+�qbp@�!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī:f����p=�3Yj>��N��x]-6j�"Hs�MH�w^����@V�RY8�,�;��/�� �-�b�+�