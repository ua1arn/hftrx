��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"��ցY$݂~o���*��b�<�Qq�T/��gaȚ�``�+c>�%�o)�[g�Y1��̒����4m����_��V?�g#A׃��45��R� \��W�Vh��=]u[��[s���;	���җ�ɸ6�����/R�����/�d�U���LK����,[����r��1��4����K��g�V}D�B�&��8y���� 0��Pxc9�\��o��Vٶ\�dD:���{�e��1ܝH[�*��I�]��
3��������ɠ�J�@Po؆���Q;��5��x�"��g"\���ĥϗ�4��ɖ
�x�	q� �a#�E5�oM`yZ�f�Y?�����G�%��N퐐��V6UF���.�bˡ5ʾl��IB������s��
��V���m�̿��Ґ�-]i���>��bq uH+�@�a�GW�+��S9d�J�aI>ʤ%��r`<�[}�I�
�}���2ݦ~��d�׎�!\:����ʇ��\���@����!�zKl��K��搑iؠ���u֦�K�q6� �kc�D�>��#�F��k-�$!z��@��Epٿ������,W�g�o���M�жLw�н%hl���2*������d?��>׈r�ዑ�ۜ�)2�_�ART����&k,�+Q��Uq��|{M-ٝ4X���0��Ml�)�+����h�xw1uux5N��r��b#��[�\C{���7z7��PGn�����7�Z��<F�)��x�4
�i>X���Z�n:�D���Z��8��~H�}�*"'@�D̥e��tX<�4?�p�<e��m�8��V�%�3�=hҞh�猿|l-x��揮U?1yB��jɩ�&�����Y�Y�]5Ŧ��kg�9��"��_�ۭ�ɕ�L(G% <���|e��W[N��"e��~�v	!F����?�7H�E������RoV��&��t�w���dDA<��� ���K�qս�GL�4k�R6˘"f~1����<="̋.F�W�8v��$�f�GQmG�M^�v��:�]{b~28�t�A���Z�����	H_�Jf�E�?�̭��ʋ�hMR:�I{�=�}l�t�>.8�x�>ס��\������@_�D"`#	S;:�ũ�٦%i(t[6�%�����֚-p:�32�+6Q6����ȋm�w7Yնdƿ������7����"͠�����`$Ź@��Ĭ��Ԁ���<�?v�I��d�j7����e�@�b�=s4��Q[g��$��g�����*,aM6�.��s�
���\����>�G�����O~�y����I�,ʣ�a��b��ǈ/��o�6�sL�&�ɖ�י�~���bw�s�ȅa3�����g�C��c�`��nW���2���W�<>�.~L���[Ϋ�,@��~J�i�Lo@��CD1e8#��i��c"���+a��@����WyB���ST�'��T����	$4���jr��wٴk|~ʪi9
���X��J��� x�?��'χ3�s�7����w�@G����v{#1��η��o�X�5D���7�߬b�A����sخ�e�M�Z1Q&/Ԩ�W^05Z,�j�(t8eI_S�gm��>]��g.']�5��g��^�jH�)_Z��l�>�_�G��C�a��_VB�{��C��4�!{�g*�7i� �f5t/s[��ȉ(%�5��ՅZHX�9b|P�Ŋ�'�;G$n�EVd�4T�C�X ���h��`�O��x�-ـ*\N+N3�o|@ӣ����j�����tԿ�f��4�k�2��-
ז=�6 y�� �ľvK݈���҉��L��Nn��`y�^�_Lu���n��4���UQ��`�al���;�po�v,�`"ʣ�@�g�����Hf���wf,���%���Z���q����0eT��(2
��UX��pݖ��,�`�B+µ�暡߫+�� ���G�ޙ|�#K������\6���&|u`�c�qv��9���V��U�2��@�Th����;��o<+ԝ���q�V�?jy��3���A_O��u�墋xƚ�d�������k��抪z4��n�!��n؃Uֵ����O�/,�P���Z�џ�1��#=c�D[�"h)l�x�h�}L{����F�h>l 
��1_�&����Q�(����؎�Y�������B��$�V:M~�T*sF 5��9"��ܸ��u��B���ڭ�(sZ�����!]ɆS�j-�Qj�`��$����%׈o\�࿌=2�F�r�^�;��*]۱��d蓨$B�F�̠���ջ:(\l�5&�Ǔ��/Y(q�>'��C/B! _�:��3�S��Fڟ�$�^�� &��K�=X�����	=3�p����e.�`$*ԏ{d�8g��}M5*�V,{q��7bO���$>d��R�1pT�Z��HI��л�N�b'T���0�ڝ�q�qPV��=��Պ������2B���CB	����7��z�ZO��hu�5��-*���l��1�~�ؚ��v@�mz�����*{�N�Bƃ&���3pH�h��c�֏����\7V����4(�B.�"/m����0�	�s�߱�n;�]��):�K
i��s��
��O�'��'���Ha�@�zjfc�j������;�M*I6f����|^��hT��(����#�-C�R젖rC�����P������:��jinB\��kQx�Z��|J��F�/J�_\�2�b�}�>kS��2d�w����^M1r����*����v76mٓ�M뮴Y�+�����8&�}VA�Xן��K:�=�g)n���ȩ���b�׈ۈ�m��Q�%�i|�,Z����a/ȳ�g2Q$�W0�?���>��Xn�ս�?-�w\�(��-]���N���Ґ�Ɏ��Z�{&�{�Pa�;��RH�M"D](�:��I�`�S�������
>./_L�;sȲ%rZ��f�d1��a����1Sӛ��\/[�P�Nr)�F	�d�e�4�.F�~Ն�����#��>���I��᡻�i%�>�A��S��� �ښݘ�#��dP
�w��F��-Ǫ)�`�N@>��[�{���Nz�fbN�!X`�-���<��2�z7��F�����n�{'�׊[�����s�>���j�C��3���$��Y��/�I�{�>V��ź~�yZC�����J�?{]PD��7F�]�������%�أ����a.ʇIK�����[:�L2��F�`9�w �4�Ӗ�7�7�	�8���[�Z���<124-*`,��`����q���2\���?*�����@�ኃ%�d�|���2؏�脊�:	r=��
�}��tRI��s�
�,J�~UIYz\N}	���Ct�30L��\'Xk�qX�4z��ԝ� ��,�+鏤����`��P���CӇ����Dݞ�,��a�X�q�_��diʨ{��y�@�1�/KI9!o���W��(gӿ���z�l-���?VE�
?ǂ�#s�<�J�o�o���b���q[���6�b�IRn?C`����|6�h�9|��Rk�n�f ��q-�#ⰰ�鷦�gҥ�Vv�C"��&~�Օk`��x�a�yL�����@(�h���OU��E=�"Q�^��7��g}�B�u����\·0E�"4��C_�)�&��;�Ru�߅TF�wW�Ӗ$�#?�%���s<�»(䑀�Ϗt@dm��=�FP���>���&7BOYrh�o�	Vboڱ���+q��Y�&]J3���_#:O�����k��\��"������к���^�,Օ=��=  \Jr����v� &Y����AO+�J�Ȍ�K̬�O���;�
�B�ٕ���?���͞�YZ�H��2�i�S��r>�t�QZwi*�p�i�P�B|'�RV�R�eR
t� n�(Mܕ��|�� @fq��	ۢ{zԇٱ�s�!;×�)JV��K5�/�>R�Gm�>~"�N'���j��
CYŻ�z1�h��Z/�-�^e��r�*�����5�	Ʌ� Fq0�	ճ�6LTc\�n����+-�e,�I�4�'Q_�p�BN�=T��uW=}� �NR���@H��%T2]����[��?��n%+E�O�!��U�?�������*�����������F@K"�n���sr>X���.���N���\^X�Q█ `b�,}�=|�� 	E\���3���t�x�o��C-�'N�a�g�)+��R��eE�g�����j�q޿.�ۖ�j"ʇ�P�;�)A�_O�6�A����.ez6cLvJ���+7�-���lQ�2�Mx��Ր��-�.f�	ٕ?pͶ?�#�G������	����"1J�����\�� >�S����'�>=���-����6����.4������9:�6�A(�GR�Y�t����[�(�ɱ������ʦ�'�^��}*�H*��E���}�e��/��?�,�d�xtcnHAGM@)�%�|ۿ�[L�\_�y�!�0�A���C��K>�E�ƞ��Eg���`f����F�tF�k)0oH����rA���_3�{#�1��d�����{ �Uy����ٶ��U��߷�Xqlfsڹ(�J�Ʊ�p.���������t_]"�4�ÆN��v$��&��[�-� �?��I�`i��xP���SD�!���66��b��,���_�<P #I�^$��FJ���J��+&{��?�'D_�4�����4M��9T@�rv\���wƜN����F3�h!C'�9?M�Z�ٚn]��QI�]�7��E����Be����^WZ�?���4�i�r���< ��f(l��"3HX}J�OԽj�����k�»k�fqur1�gY' �pu!O�u��&��i��6u8!V�Х��ᑚx������,�L�M;}j��Rլ+��6f������tm7Ev�tG���R�_��l����g�q#�(BF�@����X���<x3��J��p@Y��%-�2��C�v����?3RSjE�-,(�K��m�@S}'Eg�ƭ���"�+(5��V�ާQLp��`6|6ρ)8�:D|b'��#`3tI,�>	����;�L'>+C��{e�W0�MB�y�F	�'�����1�_#ܞP�$��ۜ/��,��y!�\]��Q�<qjJ���{e�I�ܵ1
��%�i
 ��MozJ���4�'3�9�aX"3��E��1��`'��4Jk��{j�6"L��5�C�pb�ǝ����-��ԑ�t� &��g�c�����ra8��ur�p��o�2�Ri�g5+A*ߖ��	=_g�k����eA~�л5�"-1��s�i˚��	���X�!)���첥O�� MdO~�ӡk�N���$�G>2����Mn(,ii赦�I��F����'c��jw:�W3�L��m~I���k��N��_�x��V��m�\��䔎(z� ���tS��*�ޯ�,�!�[�S��uh����	����"N�x�?�C�H�g�Z!�Gr!�)@����"��o�\��)��[�i�,��`8��+r��Gn�y��I��G�g��f�r�"<q.*�X���tw�&�'��a�q��q��N�N,D�(Y�M�v�	�eTc���i�T���+|V��}X�M��m��i�gdM�����V�?9���l(�y��g���}���D�~�D����n�A6sX�B�BOj�G��}%w^K�cp�s���9@�2�'G��5��8�P� �G�} �ǄS�])]��iM�z�s������;��j��6�O��oH���P����n��ja{��'QG,V�ϩ��wV4=_fD}��@dU��62:p�lP ޜ/�Yp���Y'�V��=��|�.�_	�3���3]#o81�s�+�Q&tze �Kx�P�mz��\D!x�i��m{E�K�u�.��U�?�6����L����Os���B��L`�o��_i�Y�i����M�0Ԏ�P����5ԙ;$H�;)F7�hέ�r���<���ab�v�!	��G���t�Y̬����']Np3p�hϒ�C���Dӭ9
���~�6�����,�ۍEw��0{1����,'2�(PUQ</L�iwYm�,����cޏ��	F�Z�[/�⾊^��~W�2�K��N%7�D>zI���y��S@�ʵ�;�lA
򰏙�{w�����r�T����*��i\7m�0��]�W|��$�f�-���s�|��[P�{g�~����J���i��q|���=�����<�W�!�nU �����Z��(����w��S�� �g�/���}b�?��x��Zӻ��qrq��RZV���l"�|�ٚt�O�*&R����S_����;���d@�s�;�撲���2����Չַ.�AQ�n�⯭�*&6���;�K[~V�w��|'0e@�D�WEq���}Ih�3�sU�y�� e�����U��շ=m����ALOT8�,����I9��Ui��<�TGCU������ ��0 �g�;���`�7��;J��"^`!��������"��@�uǉ������aL{-/�>���v1Ʃ��GO�%p-��Z8$U���"��qw��07@k�������4�N�k�X����֮�2�<)5�.���� V��e�GVRӂ���(�nJ6�����*�����`��G< t��m��V�bV��M��]�RV�*J�����e��1ub��	���Bx�ǯ�M4������uCk��7�m�^:���D�8��i(�1���Olƣ�'�����XkWӗ����y�@�_��budI,�H�b���.]���apkj-��Xt� q�m�_�f�w���=F�&��$���)RP-��t����OӴ���e�h��{�l�a�0��`Xɺ
��+��VvR �~�t��DЗ�6�<����,��)��x	1���U�չ[�o�҇��u���퐱5����r�棖G�{08\5@�9]�;6Х�{ɏ�/��`�ٚ��o:�|��`�^���9(��.5�}/�3�f؛&��SX��hE� ��/4X )�?��`�Bu��j�9��bYo(��I*7ڜ�+OnZ 7���f�=����/l..v�b|.3�ޯD�=������yv��kOC]=�P�~C8�ABy͒�$���	�#��׷�Bs�����	ޚB�U�I3{��p_�x��w���.���*���5G���
c�{�s�j5�M��XW�&���d�����S���q�dՇ�Ê-ݢ�u�X���b��`L2��K��J������͎�Л鹪a��^t�۷���co��K~��kF�A.�����[��U���}+븾|f��PSP�,qI�����7 ̵����,���z����,� �H6���-��RI�ѧ�|ϧ,7
M�{P�M�ڞu|XY��+�}	}v���k��2��T��@"�v�M�s���e1ldu"$��#�h+cB�����>�<� �Z�M�t�hJq{����i�^:8q���� 6j������2��N&����C�H�c��#5�}���q׽��MJvlcqJxK˓�P���s��[p.����H�W=E�~��n��g��%^_�%`[dX҃�+�?�w��R�+�� 1�̰ �r���r{�rp%�x��y@�DW0v�G-T��(V�tS�?��vkP��)x�l�Q"��S�T��hq���(_C��hf�ڞ���u����5�0�_��j=������">p�6p�ܚ�y�xհ�Aގ�kF�ѧ@�S��_�u(ɡ��«���QV
���v�N%Gš�,�w�J��RG�C��RJ�d�)v7����:H-��u:����S��~�mY�f�����Ϳ�3��0��ȷ �i���i_ް7޵>����HC9�(��'��D5%}��ha�+��99�5L%�CKfm��lP��y�����U��y�5���r>Vph��܋�Nm;C�Ȋ��g������7�Jn{Sg�A����<�:�j"�|��){͘��8@�6���N��$ͳR촭Ζ�_o���x�X~\������������n��mW����z�.�'P'��~s�O�9��,��!}��0@s��bTn����^[q�H��x���:U^]��(�v�oQ�j	�YA��d�g"۶��s-�r���Q<V�vڞ2�
;$Q;�9T����A#!��M,����xc��t/�4�����:M�ϧ���&�Y���5��������'߼�K�ޤ#�1�(���	P��W�{����5�Q��]p��5>�t�T���oĒ�=Җ��P��xίq&=��ϐ��Of�ՄԽ�-��y33���Jg���D.�d��|^�/�H�~]�]��㺜8$Vbr���!n�1'X�(9���u�c!=�}-��@�k�,w���7X���J�A$����L���P��Ow�*�Vu|��;��1���Φ����!���(�F���Yr��S�c�z\U~
���Q�N4��%�Ha��������͂�P�F��G�y�3h��^�4�WV7T-��\�/
�Ӈ�3:#��a�TM���]�֥~��:�3����d����+Z����U���ZV�'t�I�����i�Ð:<��[-����>�H�}�n���NZ7�����NŜ?�
ێ^�:d�Qo5�Gu>�j�w_�jq�v|��>X1�(P���xY+=驙s�3��S�Q8�j͉T�$�,(�!�\[�[�bפ�p��2e��<k��������.��Vb����;?{/i�D��¡��y�A���\�.��Q׭�"&�l��H'�ISX=wϢ�T���I��*��Ql,���$��D��.V�*�z��9 c���։�W�����Y��b�;ЖG�X�X�=3���N��z睎fC����Ϊ�]�/��7����y�P�d�|1}؆�m-�\�)�HV��V�>����6�&�^�O�9�r����_oF �ą�U��:4��u)esW�gsd��sR	�_�Y�N���퍰��{�����＠�Y+�`8J9�-VvqG���rD�WT���^�.�c&�H$fl2��I`D`����;T`��?�nȋKDj2J�U�[eN��/��u�؟ùV����۸}QZu;�����nU4!k:�@<O�Y�� ���!�����M���t�6+7	͝�x�̸N?"?�y��_G�\ߚ��;�,�_oE�x/���0���!Ni���Z�����K�8l��Q$ْ1
��M0�W�S��}��-��ݛ�T�JNA+�!���ڝ�!�x�֭�feV>�[+����>]vq]L�N8�,c�,z&8���e�@�tf��A�������բ�t��Ƕ��_�f�f�NoV����	�X�5���������q0�d_����ԭ�|,�P.1FOq��� �lD�c�E6� ��#y�1$��k��Rc1�!�_"���?*�L|/���_QUR)ٽ�a���h �e��$�/�27�@ʮ�k�D��5�8$�y�"`S��!nPI*�m9�Z�Z?��2�:���x����G^n�XJ�	Lj��H�𾓋�z6�����U�̜�����u�j�!�TJ�>Ϟ�:���6(�ס���iTL
��-.��U<"ʎr�QY��4o��M��d�;츥���x\�U:�^k��D��^���P�w�:��� ̉�2�!hٖMޠW�y^�:/�SZ�jB�f)+\�߼�F���9����&h2�2@��[.	i����B ˓���Alf�ˁ��zP����-�x⊋=���,���e�{�CQvA��k��?.%~���p�e2
���V];�_0�|	�B��
���V$�<ɿh�"p���5�g��@ۙ��=�������GCյ�`2�}`[�\¡c����uX�G����S��BZ��>�J��Ju�&����_s��P�"&.�/�Z�,�;[t #Id��#pǺ���Y���GEGK�{���}�r丕�%���|�[BL �q~Ę������y�)�O�ug��T26����ӓ��r!�٥��7�P��΢��sĜj��"ٚ�#K*`��!�F	#�ȕ�$%�OA�֌�CBo���c�
�ƹ���8��f�}~+�L΢1��\�&�B3����y�����z���2Ю�9D�u�k�C��u��}������+A���1A�Cg�vU�;q�Ϗ/o��PC*K�kf/;�XE]i���a`x(XZ�F�\��UC�ǯ_�� ��m�z2��(�� ����Q�&�0�ۜr����Uq��Cz>L+�_az8?L���(�cM��y�0kFn��Ĵ7~�h�p5�^(2	��( r-�T�j����M����NL'��ڗ��F[cg��4��c�݆���^h�c�E	6:��
����#v��������K��.�����<����Q,�HD��tlnH�;k����G�l�=�m԰�]F�֕�7�b��/���'�F����.������Cc2u5J|��T�l��i/c���~ע�'��F�4,��9���[S=y?���V����0����r��S#�l�˶��ֹ�=���O��M�6<�V-A�-K��x���Dj̀������E���jQv��ř��,0�Q�\�z�A��c̊ ���Q`c{:����jQ����㮟'���$>
ŋ[!��V_��k�JVU��Vm�:��?Edg
����)磀�n����� {�!�{#.���w|�4��i;Ы���������NY]��B.B�	��C�-_5�u��|�kQWT\���p��o��B��T0TYg����'���F���	����LR��0���[?#��ɯ5��Bů�﭂qނ9,��0ۼ����HPB(��0>�vJ�����G@���� {� �r�%��n��G�e$P�Zn'� "j�Y0�>k+J�g)\�K���ͦ��6��]�o.�u��6s^l�k�{5�p�)Nʲ�q<=ŵR�Jk�Sm-9<��_��77p�%F�%�ȧt2	Q�n0�i�nR���.d�o���&@��0P>�)ٹ��U�GI&�u`����kW���Tu(����ۍR����,��z��:@y�2� �=6��<� ��Q��tW7 ����7Zf��'�kap�DF��Ho�~i5�T��K����e�l���ת�p��8y�uZH/o��}��TU-�� ����_@�֠�Q�����m��tDb��{��K�I�dN����	<L��&c?:����"3ѹ$�Fl��UB���haz����ZET�^�_z�IK!�@�θ������@~�t")1*c G�� a��X�������ń\��.��ʇ��Y�y���"޴�F���5<��:�� k�G��� 'R�1�PxԴ��RԩCJ( ���&�RfY� 1���x�x�
� ��ᨢ>���Y+� "�}}rX�f|�̫k��dAY�*ֹ�+ �a�7�\�w|�N��S=���T'Iٚ��J_���eOƋ�$�A�m�@xB�@B�@I���Jl{o�vEV��o�K��[Es��RҮM����sP�7��ȶa�ʉ��0���^�I�r�yl���l�a ���ˠ�2 l�,5,��u!��:��_�Iߎ	460Nz(bl�{/��]�x�4�� r]����|,7�H����:i��*D�{'�}Ձ)�w��-�)_��>=Qٱ#�Mfwc�8	��BNJ8�L��i1=qj���<BUs�H�0�� �P%��ss���RH�r�~{1ǻ2�[3�Fh� �� GbbU�@±�,}w
���M�:�ā��A��ٜa�U5��Q/[�z'�����5��1;�~S;),���y�*w�T���?��j6j��ێ3&{�*��B�IS0���E����L]ҝ� h*G�(��_ӥhY[A��tGvv��!�&Z�����R���e�v�c��#�zS65��!�v�`e�?����6l�����������_��#�C��$B{j���E_�_6�
�]%�ͩ��md"˞z��Gx1b�s4�ʢۋ���ұP�8�����l%W`�HƙB���`�w�M�s�8�gr�1`a�v�É��I�b$s�x��P�a`G�1���1+��m�t�����7PJ�]��Gv��(������\T;<g�����s"b/�o���f���|v�M[��w��"���G��ս@�R�'0�J^�0]���C)#T1�P?�0����eu5M�[B2Io��s�YΪ�@��Ő�C	nM�ud|���]�O=�G=�2�+}w���F�	�	��a^����;	j���x:��rn<�.;��6 O��?�N��5^8�^�|�j�t�7ܖ��~,d��6����U�������F=���QQ�,�z�@�9C9��Nβ�iT�L\)�w;���Ih�L��1�}�o'��Ӏ���/K��)�zb�"X�����Ry��K�4���l�?upM}(��a|m���e�P�܇�S�!�x}F�Q[�olΈG�!Ʌ[N�4����|dᯒ0=RAi\�F��
]0��p/}�8�'����ĥp�P�Q��
M�d�ɜ��o��Z�FB3'�e����A�ß"�A�3��|�}�ӱ�b�Ky]� :.#FiU4(I���%�~�,r<r�Lb��v^K�Y��M��ars{�
:n�ԣ��P�z	���&�ʗL�+%�Vm��(� �9��
g�GdB^����X�Yc�T<ǃa`�����&�H|f:��.RD�݌~�\�9�}��B�B��	�"N|��׺{x�YD��'�aO��;���q����E�Y��az��4��T"+�ϓ������/��̮({Wj8mf��@���3��!�l��
�!�R��lI��'�Mr�w�g�z�f[�A�=1����L���'����/D%�X ��82�U3<T<��t�т��K�S�{��j��}2�!�e���Ą���}�8�G[o�!-�~ܪw��{-�d�ܻ��tGjL�p(��-�
�b[�h�{�լ��W�:���._�ΔL�8����7�%z���h�"9g	���.��!h�h�K_�H��_�Ύ�^��
(�O��B�B��b<��:�0�L�5���xf�V��uZ���HN��r<�W徻�(��V���瞟�܍s��9�p��N��� lV������\9oЭ�n�-��[Ԑ.|CF;ZV_<躙���Ֆd�z��1<�9iz9�-w���3[j�{����oR�V�5_@�o�A,P�nH�A��L�?�:�T���Q�؛2u�Q�]��0��AUfl��yC��j���b'��j�A��4�oE�zvG��:�;1�%�E�b�jE�0G��*�AQ.�@Zw��@;�+�p�#	�_����kH英U����u�z���m�)�_O����8;&��@P��9�c��W hjs	�פޚ��V�������#��Duj9=^Ȃ^�'�ά�؈=7.�($�"\����&������#�,RX^�i��v���U����h��7GVs�laI�ePZ+֤.�ˆ�[�ц��a�[u�v6�p�����Ϝc�
�`+�l���.I����{V�KT��Q&F���^�9������`18��u�� ��@�T�cVTx#@*�J���OƬ4��ߧ��;E!Lۄ���;܋���NO��!�\�i��Y>L�� 1ݎ��S��H�5A�2����8|9�J9�8���q�K���������@���>g�ѹU�&�:�:��T�K���jF}x��0���B��ٹ�W{�j�#�B��G:6��a�������Z���#�y_w���WO��c9�D�Hwfe�CϿ��	C0X��(��,l�X��g.���˵� I�RK��9������im�	I��v҅ ���������|���J����u���mF&F��&���펵���/�e��h��A�(�:��"�7�РH3����O>��t@�~�Sɍ�,Gx���Ϟ1I_�k���\� ��;��<��@J���U�>DY��A�F2?��\�4�B*NiU|k[}P�����{��s�I!XF�S�L�z��<�nx:�Ȥ��'�0�DF����re銥����K�{���܄f=�`�.�KWօ���4�M|���x�A;��<�5l�+ۢ�`��k��L@�V[0
��O�*�fB�8�>�|����
r�V�y�Q|6R�:X�?�YdLjo�2�3�2�7��`���v����3f&�\܈V��D�� ��eC�1�AI]/옏)�a�i��B^}^���W�3�_����7A�ͼ�6�|���Z?��g;u��[�و�M�=�R�]+:�c��=��:!w�*���۠
�:n���� ���l�}�c�/����~��,j�\�����W�"t`˒}�Y'z3>�YE�0�9�}<��  �|<�߬f0���ւ��{��IJ&�
2=��4������0�}����
>����\m1hm,&���M>ƃ�d�˳���1�C�J���g������K�K�����کS�m��!Z�@R�����o�l~F㚒W���	�q}tw.0n��y���"Z�{T�.�.��B|�$kg\��G,#�MS��2p&�%���nu-]�-�;��LwH:
C:�/u	+5;����[8\T���_z�BG��_�:�k�����5Ty.K��>\�R69���0���_	W�����O���|@��^���ǞhLXK�������<��{���[���Cơ����B)'.���5JxKی���AO)8�A��?�B�tL��v9��v9�5��j���0=��F���2�n���Fw��"�r-�g��aBl�(��t>�[���'���>�bS�W�ԟ۠�E�z�iR4Vˀ�G����@f/�\T}�Ks��.�����4W�
bʛ����Z�
�HJX*-��W�{�Uu��@I�Vv��l8[,��Pe���!�Ӭ��D��(�����-n`Ϻ�LH�?��KF��2��)���o��q�P*�����qC�s����=F�aE❤�,;�?��w.}�;!�*?�sb�)�wtd���]����l��ARm�<���X����U\�9! ��H�ε��B���w��=q��d��W�������ٱC�����FW*�w���ǘ@3:�d˴�>ig}���2���)���[�y����I�s9m��֘Ib�I|$���(Tg��UnQ�"<7�Wq��|�c[1��eL.T�T���F�������PM<7$�A��M_`��x�,�$C�G��N5�q�Br[)�^W���QJ�N�=�������Z����E��vې/ůM�!�Z[g3�ߝS�*(I��M�֨��;_��_
K�v�t�k���T�[)T@y��֖䚐��BƺD�oz��Ț�#��m�H�A�+"5��s�X�HrN��
�/.
>���t�$@�3��Қ<7�Fs;0E�wLGTB]�"�w��ɦ��C$ͮ� ���m���0{���2�1Br�m5�d��`kiA��i�`�,z�����^�K�=�_R�%v��W���?�@�"�}�V	��Pj�L���W<�f��.�2hWe����}7���oaT�B����2UB������D�a�P0��/����B��Y���a�a�,�6��J�����,ϼӣA�K�(��n���t��BC2_�t�S1�d�I�	�_p��{�B�3g�eN+���1�+F$��kO��Rm���v�L��8��~�#����S&p�D�8P� ��;�R�qh��f_�ً�_;�����"dL$�aKM�\�fC ���<�*��G�Tl���Ѐ��2X������U�f�yw���+�f\�q��Y1��NFo����	������<2s�<�� ҏ�%���!	$�[�e���w����dLĪ����My��[���8%�H~�� �TQ�Y"��s�Ez7 @.�t���aw F �c�1��4_!] �ט[�jٹt�2c�����P$��S�@?ͤ")x�g\�����Ȩ�-_��;K�˷�<�2b��2�Qp����m?�a��������c��kk�y~�.z t�9H�"Z7�a�������0)��������:��.��V�����_Re+/��Y�P���b�7��V|I����̴f$;�LCBm��9`��xzF|�juZܘ[���h�ݺ����2�ue�FN�9֫��̓��q��:�_˝ѣWE�IW����
l3�>��8`��
����~��.�6>�I'4���rsY����@�����"Cf�w̀�7ǧ��C�!�D�u�<�BXOf�&���K����t�������A�?2m͇�[���n1w��{U����q��Hl`s5ÏΓ�М�h�۞Ԟ66ɧ��S�6n�����m��d^�}�(X�:NT�����LyT������:�~�9Ds�O4����f�-�)6��<��`>�8E'��{�������0E^�Wx(\�'��ǻ�2�~5Yr@UHLi�
b0L�2����¤s�!j�z�\'�5�$0,_G�;�А�	@:i�w��4���(��{R����|~�Zc����[�0 �Ƀ
�+J8O��VC7�]<��c�)��v��P`�]eU@_d�C��(���ZG���Ļ�����ͯ�[�4M�c
F�@��q�tcޏ�`O�Ĩv��œl �$�d%�3[�&*_pf�<��z۫4
B�.Apk��4�-`*Ƨ�z�K�P�k�~34�M�����]pEzHȞ��}�S@�!n��IN�{��'�*�3R!�А�U�Y��u4���������*�j}6��R�!�?�n�����w�����s{�	����Q���=��1��� �Z�$��l���y���WYPjݤ���P���Ŗ��ܶ��6����~�s�S^�WQ���ch6^�5����=�sN"Q��6f6�F��oi���\�S�*�st�6h�wמ���t� 4ķF�����]#9��F����T��Q�b��?8��qIe1Uʕ�=��"X��<`���^���:A|˒� N����a���'�W�;���=�3�kX���d$GW�i�O�Ⱥ�٧��+�g�&Qy8ث?򣥚8-��� s�љ��0Q�P�p-�v�%1ڡQ���eY-��_��+�^i]���9F|��S�'!��n������D��?د��:&�>���M�-ԨLI�l+����G+{�
���]���/�(\:,*��b�*�÷�JV\p���{�t`���(���`�Q�L�� �UaI-3:��<q�f뱑t���l��9%�Jn�aX�x'����WQ�fL��#��"�<v����~����D}>N	�:kӷ}4r5��]K�p�]?��r��]̰�o�����,k �Vs5<�`d\-��-���ӳ6?�c=�F�}�֋��a��B_=��<\F5�f8*54=`j��Vw[L4�����2�j_dq�m˝�,���~xγ?�͑�j>��J�d `�\�!m��l�\#��� DK�����p;�W�њ����>����W1@��)K�\�>-j��ga������ղ��V��s5m�1?��u���t��l��N�*cZ����O��A[��~9T�4t<X�ec5�{7��G�r�NG�Q�[�\�*�/0���T���v�8M,la[&l��1#�MYx
��8w��_��0� ���8<�i7��b1��T橺 ?�H�h���aD��G�j� �o�Y��b��s�f��_�(���	W�iÏO6�S� �{\O�M���D��6ZO�eH�H�y��Vjw������~4��76Dk��D�MB��"͒ۯ���q	!��a	�#s�I5���$�%=�ٳ:O۸1H�3&�2WZ�C�WAv�!��^�&l�-���=H�,�^��/�0�C�X�)���tb|�;wራ����dI�Uɝ� l��諉�p��4|�����VC�.a�KP�`Ggՠ���V<��
��,������'�E�����Xc"Gb�~��ݿ���G�*����G�8�z�艒�����1��&�b��?k���<gk�aO^�{�@��5(�:����a���[O�L�"n'w`f�D�:�$�4��m䒀s�T��mvJ�����؏�X������1z�'g�|�����$k M�Ǥ;��u������$=�_�K��{���͠00���P�G5MI`�� �h�1498ۨ]��pD�^�?8��Gn�4�~Mߝ��&L�w����+���T:�}���ѿ- ݡ���%�wei�4���I�츔y8ؘ-^阯�r'����5:[}�χ_?J�z��7o���S�-텙���f�C�2!T.�!^��Q�L������\^�@J�wdmjq��+M8mI�~��(���X=�ES�!dT ]n�'A-�XJ��*i�Gm�f�,V&��w���q�ۺϵ�Id�%.b�u���[ssM)'��O���Ib'�A�2V;o��s�w:H����(�ڄ�O9��F���h'($��L��5j,ў"A�O����%��XÊ#���4,۹��I��ny�U�s<�.�`����̢-��m��L�0H%� �[���o} l��(�p~�ʡ�v=��cU߫�&V]u^, �J�`�GH��̬lZ�/�*��zO��s�t	Wf�Us��9.���UK����u��L�O����R�� �iKH����t�pvoF�����`���^>��SQW�>�؛�����W&������kf�P��U��w�z^�.��Y�q/a��Q�!�s�a=OF����?�#�o�U��!M�S��6>,X��u���
�0�YӢ����,��p�_��ӝ����8�ď�龬�Q�g~�2=m|���ʵ
�R�1g��POX`M�+&`���{ێ%	X�z��Z�n�L;/=��n�.E�x�Ќ���ȍ
K9mzC	|�")�\�_�1�zmǋ��^�8c�~.zPH
1W�9����N u"v�D�#&=�
�q�Q�`O���]�u���sr�鞘��u g��q'p>F�'|��lw%N���i~+�L�mY���rS�2���:�05cߠp{`��Z���v�sG�� aWo@3
�^��`�~��; _q�"#\	�%NIi�ﳟ�Dq��`�8����jC"�t�4���fgN������t�W(1[?��������ڻ��[A,�@tqM'��nu��8�w����-DI�Wj�o���j�-�(z\(�]+m��k#�ݲ���K>߅��a�{h���f�)�Ň(�κdn�"��LCa��-�˲�`��@��.ڙU����g2�J�]��tK�$�J�3^��p��j���A)S�+I�*I�l�Y�Sw�!Y{�il��g���V�d���J��P T�ϳͮ���Q! �aw�U>=7"=w.G�������3�-��#ѳ)��%�b�������v;9���zNY�@]�1���)����"ުw40p��k�s�|���k��UL,�`�Z�PV�(�GW&�g~:�